magic
tech gf180mcuD
magscale 1 10
timestamp 1702138369
<< metal1 >>
rect 50418 77198 50430 77250
rect 50482 77247 50494 77250
rect 51202 77247 51214 77250
rect 50482 77201 51214 77247
rect 50482 77198 50494 77201
rect 51202 77198 51214 77201
rect 51266 77198 51278 77250
rect 49746 76974 49758 77026
rect 49810 77023 49822 77026
rect 50306 77023 50318 77026
rect 49810 76977 50318 77023
rect 49810 76974 49822 76977
rect 50306 76974 50318 76977
rect 50370 76974 50382 77026
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 25790 76690 25842 76702
rect 25790 76626 25842 76638
rect 30494 76690 30546 76702
rect 30494 76626 30546 76638
rect 34526 76690 34578 76702
rect 34526 76626 34578 76638
rect 50318 76690 50370 76702
rect 50318 76626 50370 76638
rect 51214 76690 51266 76702
rect 51214 76626 51266 76638
rect 58046 76690 58098 76702
rect 58046 76626 58098 76638
rect 58830 76690 58882 76702
rect 58830 76626 58882 76638
rect 59390 76690 59442 76702
rect 59390 76626 59442 76638
rect 60062 76690 60114 76702
rect 60062 76626 60114 76638
rect 60734 76690 60786 76702
rect 60734 76626 60786 76638
rect 49970 76414 49982 76466
rect 50034 76414 50046 76466
rect 35198 76354 35250 76366
rect 35198 76290 35250 76302
rect 35982 76354 36034 76366
rect 35982 76290 36034 76302
rect 47630 76354 47682 76366
rect 47630 76290 47682 76302
rect 56702 76354 56754 76366
rect 56702 76290 56754 76302
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 50206 75682 50258 75694
rect 50206 75618 50258 75630
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 78206 64594 78258 64606
rect 78206 64530 78258 64542
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 78206 60562 78258 60574
rect 78206 60498 78258 60510
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 78206 59890 78258 59902
rect 78206 59826 78258 59838
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 78206 58210 78258 58222
rect 78206 58146 78258 58158
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 78206 50370 78258 50382
rect 78206 50306 78258 50318
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 47842 49086 47854 49138
rect 47906 49086 47918 49138
rect 44930 48974 44942 49026
rect 44994 48974 45006 49026
rect 45602 48862 45614 48914
rect 45666 48862 45678 48914
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 45614 48466 45666 48478
rect 45614 48402 45666 48414
rect 47630 48466 47682 48478
rect 47630 48402 47682 48414
rect 48750 48466 48802 48478
rect 48750 48402 48802 48414
rect 45838 48354 45890 48366
rect 45838 48290 45890 48302
rect 47742 48354 47794 48366
rect 47742 48290 47794 48302
rect 45950 48242 46002 48254
rect 45950 48178 46002 48190
rect 47406 48242 47458 48254
rect 49086 48242 49138 48254
rect 48178 48190 48190 48242
rect 48242 48190 48254 48242
rect 50866 48190 50878 48242
rect 50930 48190 50942 48242
rect 75618 48190 75630 48242
rect 75682 48190 75694 48242
rect 47406 48178 47458 48190
rect 49086 48178 49138 48190
rect 47518 48130 47570 48142
rect 47518 48066 47570 48078
rect 49534 48130 49586 48142
rect 49534 48066 49586 48078
rect 49982 48130 50034 48142
rect 49982 48066 50034 48078
rect 50542 48130 50594 48142
rect 75406 48130 75458 48142
rect 51538 48078 51550 48130
rect 51602 48078 51614 48130
rect 53666 48078 53678 48130
rect 53730 48078 53742 48130
rect 50542 48066 50594 48078
rect 75406 48066 75458 48078
rect 49422 48018 49474 48030
rect 49422 47954 49474 47966
rect 77982 48018 78034 48030
rect 77982 47954 78034 47966
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 51550 47570 51602 47582
rect 35858 47518 35870 47570
rect 35922 47518 35934 47570
rect 51550 47506 51602 47518
rect 46398 47458 46450 47470
rect 32946 47406 32958 47458
rect 33010 47406 33022 47458
rect 46398 47394 46450 47406
rect 46734 47458 46786 47470
rect 46734 47394 46786 47406
rect 47854 47458 47906 47470
rect 47854 47394 47906 47406
rect 48078 47458 48130 47470
rect 48974 47458 49026 47470
rect 49422 47458 49474 47470
rect 48290 47406 48302 47458
rect 48354 47406 48366 47458
rect 48850 47406 48862 47458
rect 48914 47406 48926 47458
rect 49186 47406 49198 47458
rect 49250 47406 49262 47458
rect 48078 47394 48130 47406
rect 48974 47394 49026 47406
rect 49422 47394 49474 47406
rect 50206 47458 50258 47470
rect 50206 47394 50258 47406
rect 51886 47458 51938 47470
rect 51886 47394 51938 47406
rect 52782 47458 52834 47470
rect 52782 47394 52834 47406
rect 30606 47346 30658 47358
rect 45502 47346 45554 47358
rect 33730 47294 33742 47346
rect 33794 47294 33806 47346
rect 30606 47282 30658 47294
rect 45502 47282 45554 47294
rect 46286 47346 46338 47358
rect 47742 47346 47794 47358
rect 47058 47294 47070 47346
rect 47122 47294 47134 47346
rect 46286 47282 46338 47294
rect 47742 47282 47794 47294
rect 49870 47346 49922 47358
rect 49870 47282 49922 47294
rect 51438 47346 51490 47358
rect 51438 47282 51490 47294
rect 51774 47346 51826 47358
rect 51774 47282 51826 47294
rect 52670 47346 52722 47358
rect 52670 47282 52722 47294
rect 53342 47346 53394 47358
rect 77858 47294 77870 47346
rect 77922 47294 77934 47346
rect 53342 47282 53394 47294
rect 30382 47234 30434 47246
rect 30382 47170 30434 47182
rect 30494 47234 30546 47246
rect 30494 47170 30546 47182
rect 45614 47234 45666 47246
rect 45614 47170 45666 47182
rect 46622 47234 46674 47246
rect 46622 47170 46674 47182
rect 47406 47234 47458 47246
rect 47406 47170 47458 47182
rect 48638 47234 48690 47246
rect 48638 47170 48690 47182
rect 49982 47234 50034 47246
rect 49982 47170 50034 47182
rect 50542 47234 50594 47246
rect 50542 47170 50594 47182
rect 77646 47234 77698 47246
rect 77646 47170 77698 47182
rect 78206 47234 78258 47246
rect 78206 47170 78258 47182
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 34526 46898 34578 46910
rect 34526 46834 34578 46846
rect 34638 46898 34690 46910
rect 34638 46834 34690 46846
rect 46622 46898 46674 46910
rect 46622 46834 46674 46846
rect 50206 46898 50258 46910
rect 50206 46834 50258 46846
rect 51102 46898 51154 46910
rect 51102 46834 51154 46846
rect 46846 46786 46898 46798
rect 29138 46734 29150 46786
rect 29202 46734 29214 46786
rect 46846 46722 46898 46734
rect 48190 46786 48242 46798
rect 48190 46722 48242 46734
rect 48302 46786 48354 46798
rect 48302 46722 48354 46734
rect 49086 46786 49138 46798
rect 49646 46786 49698 46798
rect 49410 46734 49422 46786
rect 49474 46734 49486 46786
rect 49086 46722 49138 46734
rect 49646 46722 49698 46734
rect 50094 46786 50146 46798
rect 50094 46722 50146 46734
rect 50318 46786 50370 46798
rect 50318 46722 50370 46734
rect 78206 46786 78258 46798
rect 78206 46722 78258 46734
rect 31614 46674 31666 46686
rect 28466 46622 28478 46674
rect 28530 46622 28542 46674
rect 31614 46610 31666 46622
rect 31950 46674 32002 46686
rect 31950 46610 32002 46622
rect 32286 46674 32338 46686
rect 46398 46674 46450 46686
rect 33618 46622 33630 46674
rect 33682 46622 33694 46674
rect 38322 46622 38334 46674
rect 38386 46622 38398 46674
rect 42242 46622 42254 46674
rect 42306 46622 42318 46674
rect 46162 46622 46174 46674
rect 46226 46622 46238 46674
rect 32286 46610 32338 46622
rect 46398 46610 46450 46622
rect 47630 46674 47682 46686
rect 47630 46610 47682 46622
rect 47742 46674 47794 46686
rect 47742 46610 47794 46622
rect 47966 46674 48018 46686
rect 47966 46610 48018 46622
rect 48750 46674 48802 46686
rect 50866 46622 50878 46674
rect 50930 46622 50942 46674
rect 48750 46610 48802 46622
rect 31838 46562 31890 46574
rect 34078 46562 34130 46574
rect 31266 46510 31278 46562
rect 31330 46510 31342 46562
rect 33170 46510 33182 46562
rect 33234 46510 33246 46562
rect 31838 46498 31890 46510
rect 34078 46498 34130 46510
rect 34414 46562 34466 46574
rect 46510 46562 46562 46574
rect 35522 46510 35534 46562
rect 35586 46510 35598 46562
rect 37650 46510 37662 46562
rect 37714 46510 37726 46562
rect 43026 46510 43038 46562
rect 43090 46510 43102 46562
rect 45154 46510 45166 46562
rect 45218 46510 45230 46562
rect 49746 46510 49758 46562
rect 49810 46510 49822 46562
rect 34414 46498 34466 46510
rect 46510 46498 46562 46510
rect 48862 46450 48914 46462
rect 48862 46386 48914 46398
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 37550 46114 37602 46126
rect 37550 46050 37602 46062
rect 47182 46114 47234 46126
rect 47182 46050 47234 46062
rect 47518 46114 47570 46126
rect 47518 46050 47570 46062
rect 48414 46114 48466 46126
rect 48414 46050 48466 46062
rect 33070 46002 33122 46014
rect 47630 46002 47682 46014
rect 32050 45950 32062 46002
rect 32114 45950 32126 46002
rect 41122 45950 41134 46002
rect 41186 45950 41198 46002
rect 46834 45950 46846 46002
rect 46898 45950 46910 46002
rect 33070 45938 33122 45950
rect 47630 45938 47682 45950
rect 49422 46002 49474 46014
rect 49422 45938 49474 45950
rect 51102 46002 51154 46014
rect 51102 45938 51154 45950
rect 33294 45890 33346 45902
rect 29250 45838 29262 45890
rect 29314 45838 29326 45890
rect 33294 45826 33346 45838
rect 34414 45890 34466 45902
rect 34414 45826 34466 45838
rect 34638 45890 34690 45902
rect 34638 45826 34690 45838
rect 35086 45890 35138 45902
rect 35086 45826 35138 45838
rect 35646 45890 35698 45902
rect 37214 45890 37266 45902
rect 36978 45838 36990 45890
rect 37042 45838 37054 45890
rect 35646 45826 35698 45838
rect 37214 45826 37266 45838
rect 37438 45890 37490 45902
rect 48302 45890 48354 45902
rect 38322 45838 38334 45890
rect 38386 45838 38398 45890
rect 37438 45826 37490 45838
rect 48302 45826 48354 45838
rect 48638 45890 48690 45902
rect 48638 45826 48690 45838
rect 49086 45890 49138 45902
rect 49086 45826 49138 45838
rect 50206 45890 50258 45902
rect 50206 45826 50258 45838
rect 50654 45890 50706 45902
rect 77646 45890 77698 45902
rect 51986 45838 51998 45890
rect 52050 45838 52062 45890
rect 50654 45826 50706 45838
rect 77646 45826 77698 45838
rect 35534 45778 35586 45790
rect 47966 45778 48018 45790
rect 51438 45778 51490 45790
rect 29922 45726 29934 45778
rect 29986 45726 29998 45778
rect 38994 45726 39006 45778
rect 39058 45726 39070 45778
rect 49298 45726 49310 45778
rect 49362 45726 49374 45778
rect 35534 45714 35586 45726
rect 47966 45714 48018 45726
rect 51438 45714 51490 45726
rect 77422 45778 77474 45790
rect 77422 45714 77474 45726
rect 78206 45778 78258 45790
rect 78206 45714 78258 45726
rect 35422 45666 35474 45678
rect 33618 45614 33630 45666
rect 33682 45614 33694 45666
rect 34066 45614 34078 45666
rect 34130 45614 34142 45666
rect 35422 45602 35474 45614
rect 46958 45666 47010 45678
rect 46958 45602 47010 45614
rect 48078 45666 48130 45678
rect 51550 45666 51602 45678
rect 49858 45614 49870 45666
rect 49922 45614 49934 45666
rect 48078 45602 48130 45614
rect 51550 45602 51602 45614
rect 51662 45666 51714 45678
rect 51662 45602 51714 45614
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 33294 45330 33346 45342
rect 33294 45266 33346 45278
rect 34190 45330 34242 45342
rect 34190 45266 34242 45278
rect 38782 45330 38834 45342
rect 38782 45266 38834 45278
rect 48862 45330 48914 45342
rect 48862 45266 48914 45278
rect 49422 45330 49474 45342
rect 49970 45278 49982 45330
rect 50034 45278 50046 45330
rect 49422 45266 49474 45278
rect 31614 45218 31666 45230
rect 31614 45154 31666 45166
rect 34302 45218 34354 45230
rect 46062 45218 46114 45230
rect 35298 45166 35310 45218
rect 35362 45166 35374 45218
rect 36306 45166 36318 45218
rect 36370 45166 36382 45218
rect 50194 45166 50206 45218
rect 50258 45166 50270 45218
rect 50642 45166 50654 45218
rect 50706 45166 50718 45218
rect 34302 45154 34354 45166
rect 46062 45154 46114 45166
rect 31950 45106 32002 45118
rect 33182 45106 33234 45118
rect 31042 45054 31054 45106
rect 31106 45054 31118 45106
rect 32162 45054 32174 45106
rect 32226 45054 32238 45106
rect 31950 45042 32002 45054
rect 33182 45042 33234 45054
rect 33406 45106 33458 45118
rect 33406 45042 33458 45054
rect 33630 45106 33682 45118
rect 38446 45106 38498 45118
rect 39342 45106 39394 45118
rect 45838 45106 45890 45118
rect 47070 45106 47122 45118
rect 49870 45106 49922 45118
rect 33842 45054 33854 45106
rect 33906 45054 33918 45106
rect 34738 45054 34750 45106
rect 34802 45054 34814 45106
rect 36418 45054 36430 45106
rect 36482 45054 36494 45106
rect 38882 45054 38894 45106
rect 38946 45054 38958 45106
rect 39554 45054 39566 45106
rect 39618 45054 39630 45106
rect 46386 45054 46398 45106
rect 46450 45054 46462 45106
rect 47954 45054 47966 45106
rect 48018 45054 48030 45106
rect 51426 45054 51438 45106
rect 51490 45054 51502 45106
rect 52098 45054 52110 45106
rect 52162 45054 52174 45106
rect 75618 45054 75630 45106
rect 75682 45054 75694 45106
rect 33630 45042 33682 45054
rect 38446 45042 38498 45054
rect 39342 45042 39394 45054
rect 45838 45042 45890 45054
rect 47070 45042 47122 45054
rect 49870 45042 49922 45054
rect 45950 44994 46002 45006
rect 75406 44994 75458 45006
rect 30930 44942 30942 44994
rect 30994 44942 31006 44994
rect 47842 44942 47854 44994
rect 47906 44942 47918 44994
rect 54226 44942 54238 44994
rect 54290 44942 54302 44994
rect 45950 44930 46002 44942
rect 75406 44930 75458 44942
rect 77982 44994 78034 45006
rect 77982 44930 78034 44942
rect 31726 44882 31778 44894
rect 30594 44830 30606 44882
rect 30658 44830 30670 44882
rect 31726 44818 31778 44830
rect 37886 44882 37938 44894
rect 37886 44818 37938 44830
rect 38670 44882 38722 44894
rect 38670 44818 38722 44830
rect 39230 44882 39282 44894
rect 39230 44818 39282 44830
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 35534 44546 35586 44558
rect 35534 44482 35586 44494
rect 46398 44546 46450 44558
rect 46398 44482 46450 44494
rect 49870 44546 49922 44558
rect 49870 44482 49922 44494
rect 50318 44546 50370 44558
rect 50318 44482 50370 44494
rect 51886 44546 51938 44558
rect 51886 44482 51938 44494
rect 44830 44434 44882 44446
rect 39778 44382 39790 44434
rect 39842 44382 39854 44434
rect 44258 44382 44270 44434
rect 44322 44382 44334 44434
rect 44830 44370 44882 44382
rect 51326 44434 51378 44446
rect 51326 44370 51378 44382
rect 53342 44434 53394 44446
rect 53342 44370 53394 44382
rect 34638 44322 34690 44334
rect 34638 44258 34690 44270
rect 34750 44322 34802 44334
rect 39006 44322 39058 44334
rect 35074 44270 35086 44322
rect 35138 44270 35150 44322
rect 34750 44258 34802 44270
rect 39006 44258 39058 44270
rect 39230 44322 39282 44334
rect 39230 44258 39282 44270
rect 39566 44322 39618 44334
rect 45278 44322 45330 44334
rect 39890 44270 39902 44322
rect 39954 44270 39966 44322
rect 41458 44270 41470 44322
rect 41522 44270 41534 44322
rect 39566 44258 39618 44270
rect 45278 44258 45330 44270
rect 45838 44322 45890 44334
rect 45838 44258 45890 44270
rect 46510 44322 46562 44334
rect 46510 44258 46562 44270
rect 50430 44322 50482 44334
rect 51998 44322 52050 44334
rect 51090 44270 51102 44322
rect 51154 44270 51166 44322
rect 50430 44258 50482 44270
rect 51998 44258 52050 44270
rect 34862 44210 34914 44222
rect 34862 44146 34914 44158
rect 38670 44210 38722 44222
rect 45390 44210 45442 44222
rect 42130 44158 42142 44210
rect 42194 44158 42206 44210
rect 38670 44146 38722 44158
rect 45390 44146 45442 44158
rect 45614 44210 45666 44222
rect 45614 44146 45666 44158
rect 49758 44210 49810 44222
rect 49758 44146 49810 44158
rect 51438 44210 51490 44222
rect 51438 44146 51490 44158
rect 52670 44210 52722 44222
rect 52670 44146 52722 44158
rect 52782 44210 52834 44222
rect 52782 44146 52834 44158
rect 39118 44098 39170 44110
rect 39118 44034 39170 44046
rect 44942 44098 44994 44110
rect 44942 44034 44994 44046
rect 46398 44098 46450 44110
rect 46398 44034 46450 44046
rect 50318 44098 50370 44110
rect 50318 44034 50370 44046
rect 51886 44098 51938 44110
rect 51886 44034 51938 44046
rect 53006 44098 53058 44110
rect 53006 44034 53058 44046
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 78206 43762 78258 43774
rect 78206 43698 78258 43710
rect 40238 43650 40290 43662
rect 34290 43598 34302 43650
rect 34354 43598 34366 43650
rect 40238 43586 40290 43598
rect 40350 43650 40402 43662
rect 43362 43598 43374 43650
rect 43426 43598 43438 43650
rect 40350 43586 40402 43598
rect 31054 43538 31106 43550
rect 31726 43538 31778 43550
rect 33966 43538 34018 43550
rect 31266 43486 31278 43538
rect 31330 43486 31342 43538
rect 31938 43486 31950 43538
rect 32002 43486 32014 43538
rect 31054 43474 31106 43486
rect 31726 43474 31778 43486
rect 33966 43474 34018 43486
rect 37886 43538 37938 43550
rect 37886 43474 37938 43486
rect 38446 43538 38498 43550
rect 39790 43538 39842 43550
rect 51326 43538 51378 43550
rect 39330 43486 39342 43538
rect 39394 43486 39406 43538
rect 42578 43486 42590 43538
rect 42642 43486 42654 43538
rect 38446 43474 38498 43486
rect 39790 43474 39842 43486
rect 51326 43474 51378 43486
rect 46286 43426 46338 43438
rect 45490 43374 45502 43426
rect 45554 43374 45566 43426
rect 50866 43374 50878 43426
rect 50930 43374 50942 43426
rect 46286 43362 46338 43374
rect 30718 43314 30770 43326
rect 30718 43250 30770 43262
rect 30830 43314 30882 43326
rect 30830 43250 30882 43262
rect 31614 43314 31666 43326
rect 31614 43250 31666 43262
rect 38110 43314 38162 43326
rect 38110 43250 38162 43262
rect 38558 43314 38610 43326
rect 38558 43250 38610 43262
rect 38670 43314 38722 43326
rect 38670 43250 38722 43262
rect 39566 43314 39618 43326
rect 39566 43250 39618 43262
rect 39902 43314 39954 43326
rect 39902 43250 39954 43262
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 37886 42978 37938 42990
rect 37886 42914 37938 42926
rect 47406 42978 47458 42990
rect 47406 42914 47458 42926
rect 51102 42978 51154 42990
rect 51102 42914 51154 42926
rect 51326 42978 51378 42990
rect 51326 42914 51378 42926
rect 51886 42978 51938 42990
rect 51886 42914 51938 42926
rect 52782 42978 52834 42990
rect 52782 42914 52834 42926
rect 36318 42866 36370 42878
rect 29922 42814 29934 42866
rect 29986 42814 29998 42866
rect 32050 42814 32062 42866
rect 32114 42814 32126 42866
rect 36318 42802 36370 42814
rect 37214 42866 37266 42878
rect 50542 42866 50594 42878
rect 42018 42814 42030 42866
rect 42082 42814 42094 42866
rect 37214 42802 37266 42814
rect 50542 42802 50594 42814
rect 33294 42754 33346 42766
rect 29250 42702 29262 42754
rect 29314 42702 29326 42754
rect 33294 42690 33346 42702
rect 36430 42754 36482 42766
rect 36430 42690 36482 42702
rect 37438 42754 37490 42766
rect 37438 42690 37490 42702
rect 37662 42754 37714 42766
rect 45950 42754 46002 42766
rect 38770 42702 38782 42754
rect 38834 42702 38846 42754
rect 37662 42690 37714 42702
rect 45950 42690 46002 42702
rect 46846 42754 46898 42766
rect 46846 42690 46898 42702
rect 52670 42754 52722 42766
rect 52670 42690 52722 42702
rect 33070 42642 33122 42654
rect 33070 42578 33122 42590
rect 33518 42642 33570 42654
rect 33518 42578 33570 42590
rect 33742 42642 33794 42654
rect 33742 42578 33794 42590
rect 47182 42642 47234 42654
rect 47182 42578 47234 42590
rect 50654 42642 50706 42654
rect 50654 42578 50706 42590
rect 51550 42642 51602 42654
rect 51550 42578 51602 42590
rect 51662 42642 51714 42654
rect 51662 42578 51714 42590
rect 33854 42530 33906 42542
rect 33854 42466 33906 42478
rect 38334 42530 38386 42542
rect 38334 42466 38386 42478
rect 45614 42530 45666 42542
rect 45614 42466 45666 42478
rect 46286 42530 46338 42542
rect 50430 42530 50482 42542
rect 47730 42478 47742 42530
rect 47794 42478 47806 42530
rect 46286 42466 46338 42478
rect 50430 42466 50482 42478
rect 52782 42530 52834 42542
rect 52782 42466 52834 42478
rect 53454 42530 53506 42542
rect 53454 42466 53506 42478
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 31154 42142 31166 42194
rect 31218 42142 31230 42194
rect 44594 42142 44606 42194
rect 44658 42142 44670 42194
rect 49086 42082 49138 42094
rect 51426 42030 51438 42082
rect 51490 42030 51502 42082
rect 49086 42018 49138 42030
rect 31726 41970 31778 41982
rect 39118 41970 39170 41982
rect 28018 41918 28030 41970
rect 28082 41918 28094 41970
rect 32386 41918 32398 41970
rect 32450 41918 32462 41970
rect 38546 41918 38558 41970
rect 38610 41918 38622 41970
rect 38882 41918 38894 41970
rect 38946 41918 38958 41970
rect 31726 41906 31778 41918
rect 39118 41906 39170 41918
rect 39342 41970 39394 41982
rect 39342 41906 39394 41918
rect 39566 41970 39618 41982
rect 39566 41906 39618 41918
rect 40798 41970 40850 41982
rect 40798 41906 40850 41918
rect 41134 41970 41186 41982
rect 41134 41906 41186 41918
rect 41358 41970 41410 41982
rect 41358 41906 41410 41918
rect 44942 41970 44994 41982
rect 48750 41970 48802 41982
rect 45266 41918 45278 41970
rect 45330 41918 45342 41970
rect 50642 41918 50654 41970
rect 50706 41918 50718 41970
rect 75618 41918 75630 41970
rect 75682 41918 75694 41970
rect 44942 41906 44994 41918
rect 48750 41906 48802 41918
rect 32174 41858 32226 41870
rect 41022 41858 41074 41870
rect 75294 41858 75346 41870
rect 28690 41806 28702 41858
rect 28754 41806 28766 41858
rect 30818 41806 30830 41858
rect 30882 41806 30894 41858
rect 33506 41806 33518 41858
rect 33570 41806 33582 41858
rect 46050 41806 46062 41858
rect 46114 41806 46126 41858
rect 48178 41806 48190 41858
rect 48242 41806 48254 41858
rect 53554 41806 53566 41858
rect 53618 41806 53630 41858
rect 32174 41794 32226 41806
rect 41022 41794 41074 41806
rect 75294 41794 75346 41806
rect 77982 41858 78034 41870
rect 77982 41794 78034 41806
rect 31502 41746 31554 41758
rect 31502 41682 31554 41694
rect 32062 41746 32114 41758
rect 32062 41682 32114 41694
rect 39678 41746 39730 41758
rect 39678 41682 39730 41694
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 30606 41410 30658 41422
rect 30606 41346 30658 41358
rect 30942 41410 30994 41422
rect 30942 41346 30994 41358
rect 33406 41410 33458 41422
rect 33406 41346 33458 41358
rect 38334 41410 38386 41422
rect 38334 41346 38386 41358
rect 38558 41410 38610 41422
rect 38558 41346 38610 41358
rect 38670 41410 38722 41422
rect 38670 41346 38722 41358
rect 45614 41410 45666 41422
rect 45614 41346 45666 41358
rect 45950 41410 46002 41422
rect 45950 41346 46002 41358
rect 32398 41298 32450 41310
rect 39106 41246 39118 41298
rect 39170 41246 39182 41298
rect 41234 41246 41246 41298
rect 41298 41246 41310 41298
rect 49298 41246 49310 41298
rect 49362 41246 49374 41298
rect 32398 41234 32450 41246
rect 30718 41186 30770 41198
rect 43486 41186 43538 41198
rect 31154 41134 31166 41186
rect 31218 41134 31230 41186
rect 32946 41134 32958 41186
rect 33010 41134 33022 41186
rect 37426 41134 37438 41186
rect 37490 41134 37502 41186
rect 38098 41134 38110 41186
rect 38162 41134 38174 41186
rect 42018 41134 42030 41186
rect 42082 41134 42094 41186
rect 42802 41134 42814 41186
rect 42866 41134 42878 41186
rect 44146 41134 44158 41186
rect 44210 41134 44222 41186
rect 46386 41134 46398 41186
rect 46450 41134 46462 41186
rect 30718 41122 30770 41134
rect 43486 41122 43538 41134
rect 32734 41074 32786 41086
rect 32498 41022 32510 41074
rect 32562 41022 32574 41074
rect 32734 41010 32786 41022
rect 37662 41074 37714 41086
rect 37662 41010 37714 41022
rect 43038 41074 43090 41086
rect 43038 41010 43090 41022
rect 43822 41074 43874 41086
rect 43822 41010 43874 41022
rect 45838 41074 45890 41086
rect 77646 41074 77698 41086
rect 47170 41022 47182 41074
rect 47234 41022 47246 41074
rect 45838 41010 45890 41022
rect 77646 41010 77698 41022
rect 77870 41074 77922 41086
rect 77870 41010 77922 41022
rect 78206 41074 78258 41086
rect 78206 41010 78258 41022
rect 43934 40962 43986 40974
rect 43934 40898 43986 40910
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 31726 40626 31778 40638
rect 31726 40562 31778 40574
rect 41470 40626 41522 40638
rect 46398 40626 46450 40638
rect 41682 40574 41694 40626
rect 41746 40574 41758 40626
rect 41470 40562 41522 40574
rect 46398 40562 46450 40574
rect 75294 40626 75346 40638
rect 75294 40562 75346 40574
rect 34638 40514 34690 40526
rect 42254 40514 42306 40526
rect 47966 40514 48018 40526
rect 34290 40462 34302 40514
rect 34354 40462 34366 40514
rect 37090 40462 37102 40514
rect 37154 40462 37166 40514
rect 38994 40462 39006 40514
rect 39058 40462 39070 40514
rect 43362 40462 43374 40514
rect 43426 40462 43438 40514
rect 49522 40462 49534 40514
rect 49586 40462 49598 40514
rect 77298 40462 77310 40514
rect 77362 40462 77374 40514
rect 34638 40450 34690 40462
rect 42254 40450 42306 40462
rect 47966 40450 48018 40462
rect 31614 40402 31666 40414
rect 31614 40338 31666 40350
rect 31838 40402 31890 40414
rect 31838 40338 31890 40350
rect 32174 40402 32226 40414
rect 37874 40350 37886 40402
rect 37938 40350 37950 40402
rect 39218 40350 39230 40402
rect 39282 40350 39294 40402
rect 42690 40350 42702 40402
rect 42754 40350 42766 40402
rect 47730 40350 47742 40402
rect 47794 40350 47806 40402
rect 48850 40350 48862 40402
rect 48914 40350 48926 40402
rect 75618 40350 75630 40402
rect 75682 40350 75694 40402
rect 32174 40338 32226 40350
rect 34962 40238 34974 40290
rect 35026 40238 35038 40290
rect 45490 40238 45502 40290
rect 45554 40238 45566 40290
rect 46498 40238 46510 40290
rect 46562 40238 46574 40290
rect 51650 40238 51662 40290
rect 51714 40238 51726 40290
rect 42030 40178 42082 40190
rect 42030 40114 42082 40126
rect 46174 40178 46226 40190
rect 46174 40114 46226 40126
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 30382 39842 30434 39854
rect 30382 39778 30434 39790
rect 30606 39842 30658 39854
rect 31502 39842 31554 39854
rect 32398 39842 32450 39854
rect 31154 39790 31166 39842
rect 31218 39790 31230 39842
rect 32050 39790 32062 39842
rect 32114 39790 32126 39842
rect 30606 39778 30658 39790
rect 31502 39778 31554 39790
rect 32398 39778 32450 39790
rect 32958 39842 33010 39854
rect 43586 39790 43598 39842
rect 43650 39790 43662 39842
rect 32958 39778 33010 39790
rect 33070 39730 33122 39742
rect 39330 39678 39342 39730
rect 39394 39678 39406 39730
rect 42914 39678 42926 39730
rect 42978 39678 42990 39730
rect 33070 39666 33122 39678
rect 31726 39618 31778 39630
rect 30818 39566 30830 39618
rect 30882 39566 30894 39618
rect 31726 39554 31778 39566
rect 32622 39618 32674 39630
rect 32622 39554 32674 39566
rect 35758 39618 35810 39630
rect 42130 39566 42142 39618
rect 42194 39566 42206 39618
rect 43250 39566 43262 39618
rect 43314 39566 43326 39618
rect 35758 39554 35810 39566
rect 30270 39506 30322 39518
rect 30270 39442 30322 39454
rect 33182 39506 33234 39518
rect 41458 39454 41470 39506
rect 41522 39454 41534 39506
rect 33182 39442 33234 39454
rect 35422 39394 35474 39406
rect 35422 39330 35474 39342
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 35422 39058 35474 39070
rect 35074 39006 35086 39058
rect 35138 39006 35150 39058
rect 35422 38994 35474 39006
rect 37774 39058 37826 39070
rect 37774 38994 37826 39006
rect 37102 38946 37154 38958
rect 30370 38894 30382 38946
rect 30434 38894 30446 38946
rect 37102 38882 37154 38894
rect 41134 38946 41186 38958
rect 41134 38882 41186 38894
rect 40350 38834 40402 38846
rect 29698 38782 29710 38834
rect 29762 38782 29774 38834
rect 37986 38782 37998 38834
rect 38050 38782 38062 38834
rect 39442 38782 39454 38834
rect 39506 38782 39518 38834
rect 40350 38770 40402 38782
rect 40910 38834 40962 38846
rect 40910 38770 40962 38782
rect 32498 38670 32510 38722
rect 32562 38670 32574 38722
rect 36978 38670 36990 38722
rect 37042 38670 37054 38722
rect 39778 38670 39790 38722
rect 39842 38670 39854 38722
rect 41234 38670 41246 38722
rect 41298 38670 41310 38722
rect 37326 38610 37378 38622
rect 37326 38546 37378 38558
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 35534 38274 35586 38286
rect 35534 38210 35586 38222
rect 30034 38110 30046 38162
rect 30098 38110 30110 38162
rect 31490 38110 31502 38162
rect 31554 38110 31566 38162
rect 39554 38110 39566 38162
rect 39618 38110 39630 38162
rect 35758 38050 35810 38062
rect 31602 37998 31614 38050
rect 31666 37998 31678 38050
rect 35970 37998 35982 38050
rect 36034 37998 36046 38050
rect 36978 37998 36990 38050
rect 37042 37998 37054 38050
rect 35758 37986 35810 37998
rect 30158 37938 30210 37950
rect 30158 37874 30210 37886
rect 30382 37938 30434 37950
rect 30382 37874 30434 37886
rect 30718 37938 30770 37950
rect 30718 37874 30770 37886
rect 35422 37938 35474 37950
rect 35422 37874 35474 37886
rect 36430 37826 36482 37838
rect 36430 37762 36482 37774
rect 78206 37826 78258 37838
rect 78206 37762 78258 37774
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 40350 37490 40402 37502
rect 38546 37438 38558 37490
rect 38610 37438 38622 37490
rect 40350 37426 40402 37438
rect 29698 37326 29710 37378
rect 29762 37326 29774 37378
rect 37998 37266 38050 37278
rect 29026 37214 29038 37266
rect 29090 37214 29102 37266
rect 34738 37214 34750 37266
rect 34802 37214 34814 37266
rect 37998 37202 38050 37214
rect 39454 37266 39506 37278
rect 39454 37202 39506 37214
rect 39566 37266 39618 37278
rect 39566 37202 39618 37214
rect 39678 37266 39730 37278
rect 39678 37202 39730 37214
rect 40126 37266 40178 37278
rect 40126 37202 40178 37214
rect 31826 37102 31838 37154
rect 31890 37102 31902 37154
rect 35522 37102 35534 37154
rect 35586 37102 35598 37154
rect 37650 37102 37662 37154
rect 37714 37102 37726 37154
rect 38222 37042 38274 37054
rect 38222 36978 38274 36990
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 36990 36706 37042 36718
rect 36990 36642 37042 36654
rect 37998 36706 38050 36718
rect 37998 36642 38050 36654
rect 38110 36706 38162 36718
rect 38110 36642 38162 36654
rect 38334 36706 38386 36718
rect 38334 36642 38386 36654
rect 41022 36706 41074 36718
rect 41022 36642 41074 36654
rect 38894 36594 38946 36606
rect 34290 36542 34302 36594
rect 34354 36542 34366 36594
rect 36418 36542 36430 36594
rect 36482 36542 36494 36594
rect 38894 36530 38946 36542
rect 42814 36594 42866 36606
rect 42814 36530 42866 36542
rect 32510 36482 32562 36494
rect 38446 36482 38498 36494
rect 33618 36430 33630 36482
rect 33682 36430 33694 36482
rect 32510 36418 32562 36430
rect 38446 36418 38498 36430
rect 39118 36482 39170 36494
rect 39118 36418 39170 36430
rect 39678 36482 39730 36494
rect 39678 36418 39730 36430
rect 40014 36482 40066 36494
rect 40014 36418 40066 36430
rect 40350 36482 40402 36494
rect 40350 36418 40402 36430
rect 40686 36482 40738 36494
rect 40686 36418 40738 36430
rect 41134 36482 41186 36494
rect 41134 36418 41186 36430
rect 41358 36482 41410 36494
rect 41358 36418 41410 36430
rect 41582 36482 41634 36494
rect 41794 36430 41806 36482
rect 41858 36430 41870 36482
rect 42578 36430 42590 36482
rect 42642 36430 42654 36482
rect 41582 36418 41634 36430
rect 37102 36370 37154 36382
rect 37102 36306 37154 36318
rect 37326 36370 37378 36382
rect 42926 36370 42978 36382
rect 39330 36318 39342 36370
rect 39394 36318 39406 36370
rect 37326 36306 37378 36318
rect 42926 36306 42978 36318
rect 39902 36258 39954 36270
rect 32162 36206 32174 36258
rect 32226 36206 32238 36258
rect 39902 36194 39954 36206
rect 40238 36258 40290 36270
rect 40238 36194 40290 36206
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 43250 35758 43262 35810
rect 43314 35758 43326 35810
rect 42466 35646 42478 35698
rect 42530 35646 42542 35698
rect 45378 35534 45390 35586
rect 45442 35534 45454 35586
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 42914 35086 42926 35138
rect 42978 35086 42990 35138
rect 32050 34974 32062 35026
rect 32114 34974 32126 35026
rect 41458 34974 41470 35026
rect 41522 34974 41534 35026
rect 42578 34974 42590 35026
rect 42642 34974 42654 35026
rect 29138 34862 29150 34914
rect 29202 34862 29214 34914
rect 38658 34862 38670 34914
rect 38722 34862 38734 34914
rect 42242 34862 42254 34914
rect 42306 34862 42318 34914
rect 32398 34802 32450 34814
rect 29922 34750 29934 34802
rect 29986 34750 29998 34802
rect 39330 34750 39342 34802
rect 39394 34750 39406 34802
rect 32398 34738 32450 34750
rect 32510 34690 32562 34702
rect 32510 34626 32562 34638
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 31390 34354 31442 34366
rect 31390 34290 31442 34302
rect 35422 34354 35474 34366
rect 35422 34290 35474 34302
rect 37102 34354 37154 34366
rect 37102 34290 37154 34302
rect 41246 34354 41298 34366
rect 41246 34290 41298 34302
rect 32398 34242 32450 34254
rect 32398 34178 32450 34190
rect 32510 34242 32562 34254
rect 39790 34242 39842 34254
rect 42702 34242 42754 34254
rect 35074 34190 35086 34242
rect 35138 34190 35150 34242
rect 37426 34190 37438 34242
rect 37490 34190 37502 34242
rect 40898 34190 40910 34242
rect 40962 34190 40974 34242
rect 32510 34178 32562 34190
rect 39790 34178 39842 34190
rect 42702 34178 42754 34190
rect 43262 34242 43314 34254
rect 43262 34178 43314 34190
rect 31502 34130 31554 34142
rect 39902 34130 39954 34142
rect 33394 34078 33406 34130
rect 33458 34078 33470 34130
rect 31502 34066 31554 34078
rect 39902 34066 39954 34078
rect 40238 34130 40290 34142
rect 40238 34066 40290 34078
rect 42142 34130 42194 34142
rect 42142 34066 42194 34078
rect 42366 34130 42418 34142
rect 42366 34066 42418 34078
rect 43038 34130 43090 34142
rect 43038 34066 43090 34078
rect 43150 34018 43202 34030
rect 43150 33954 43202 33966
rect 31390 33906 31442 33918
rect 31390 33842 31442 33854
rect 31726 33906 31778 33918
rect 31726 33842 31778 33854
rect 32398 33906 32450 33918
rect 32398 33842 32450 33854
rect 33630 33906 33682 33918
rect 33630 33842 33682 33854
rect 33854 33906 33906 33918
rect 33854 33842 33906 33854
rect 33966 33906 34018 33918
rect 33966 33842 34018 33854
rect 40126 33906 40178 33918
rect 41794 33854 41806 33906
rect 41858 33854 41870 33906
rect 40126 33842 40178 33854
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 33182 33570 33234 33582
rect 33182 33506 33234 33518
rect 31390 33458 31442 33470
rect 34738 33406 34750 33458
rect 34802 33406 34814 33458
rect 37426 33406 37438 33458
rect 37490 33406 37502 33458
rect 40562 33406 40574 33458
rect 40626 33406 40638 33458
rect 31390 33394 31442 33406
rect 31278 33346 31330 33358
rect 31278 33282 31330 33294
rect 32174 33346 32226 33358
rect 32722 33294 32734 33346
rect 32786 33294 32798 33346
rect 33954 33294 33966 33346
rect 34018 33294 34030 33346
rect 34962 33294 34974 33346
rect 35026 33294 35038 33346
rect 36194 33294 36206 33346
rect 36258 33294 36270 33346
rect 39218 33294 39230 33346
rect 39282 33294 39294 33346
rect 32174 33282 32226 33294
rect 31614 33234 31666 33246
rect 31614 33170 31666 33182
rect 31838 33234 31890 33246
rect 32510 33234 32562 33246
rect 37774 33234 37826 33246
rect 32274 33182 32286 33234
rect 32338 33182 32350 33234
rect 34066 33182 34078 33234
rect 34130 33182 34142 33234
rect 35634 33182 35646 33234
rect 35698 33182 35710 33234
rect 31838 33170 31890 33182
rect 32510 33170 32562 33182
rect 37774 33170 37826 33182
rect 44046 33234 44098 33246
rect 44046 33170 44098 33182
rect 37550 33122 37602 33134
rect 35970 33070 35982 33122
rect 36034 33070 36046 33122
rect 37550 33058 37602 33070
rect 43822 33122 43874 33134
rect 43822 33058 43874 33070
rect 43934 33122 43986 33134
rect 43934 33058 43986 33070
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 34626 32622 34638 32674
rect 34690 32622 34702 32674
rect 31950 32562 32002 32574
rect 30930 32510 30942 32562
rect 30994 32510 31006 32562
rect 31950 32498 32002 32510
rect 32174 32562 32226 32574
rect 39790 32562 39842 32574
rect 38322 32510 38334 32562
rect 38386 32510 38398 32562
rect 44146 32510 44158 32562
rect 44210 32510 44222 32562
rect 32174 32498 32226 32510
rect 39790 32498 39842 32510
rect 40014 32450 40066 32462
rect 31042 32398 31054 32450
rect 31106 32398 31118 32450
rect 41346 32398 41358 32450
rect 41410 32398 41422 32450
rect 43474 32398 43486 32450
rect 43538 32398 43550 32450
rect 40014 32386 40066 32398
rect 30706 32286 30718 32338
rect 30770 32286 30782 32338
rect 32498 32286 32510 32338
rect 32562 32286 32574 32338
rect 40338 32286 40350 32338
rect 40402 32286 40414 32338
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 30718 32002 30770 32014
rect 30718 31938 30770 31950
rect 39678 32002 39730 32014
rect 39678 31938 39730 31950
rect 43150 32002 43202 32014
rect 43150 31938 43202 31950
rect 45054 32002 45106 32014
rect 45054 31938 45106 31950
rect 43486 31890 43538 31902
rect 31490 31838 31502 31890
rect 31554 31838 31566 31890
rect 33618 31838 33630 31890
rect 33682 31838 33694 31890
rect 43486 31826 43538 31838
rect 43598 31890 43650 31902
rect 43598 31826 43650 31838
rect 39118 31778 39170 31790
rect 43262 31778 43314 31790
rect 34402 31726 34414 31778
rect 34466 31726 34478 31778
rect 36978 31726 36990 31778
rect 37042 31726 37054 31778
rect 37986 31726 37998 31778
rect 38050 31726 38062 31778
rect 39554 31726 39566 31778
rect 39618 31726 39630 31778
rect 42130 31726 42142 31778
rect 42194 31726 42206 31778
rect 39118 31714 39170 31726
rect 43262 31714 43314 31726
rect 44830 31778 44882 31790
rect 44830 31714 44882 31726
rect 37090 31614 37102 31666
rect 37154 31614 37166 31666
rect 38546 31614 38558 31666
rect 38610 31614 38622 31666
rect 41010 31614 41022 31666
rect 41074 31614 41086 31666
rect 42018 31614 42030 31666
rect 42082 31614 42094 31666
rect 30494 31554 30546 31566
rect 30494 31490 30546 31502
rect 30606 31554 30658 31566
rect 39006 31554 39058 31566
rect 37202 31502 37214 31554
rect 37266 31502 37278 31554
rect 45378 31502 45390 31554
rect 45442 31502 45454 31554
rect 30606 31490 30658 31502
rect 39006 31490 39058 31502
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 32398 31218 32450 31230
rect 34302 31218 34354 31230
rect 33058 31166 33070 31218
rect 33122 31166 33134 31218
rect 32398 31154 32450 31166
rect 34302 31154 34354 31166
rect 35870 31218 35922 31230
rect 35870 31154 35922 31166
rect 36094 31218 36146 31230
rect 36094 31154 36146 31166
rect 36318 31106 36370 31118
rect 28802 31054 28814 31106
rect 28866 31054 28878 31106
rect 33954 31054 33966 31106
rect 34018 31054 34030 31106
rect 37426 31054 37438 31106
rect 37490 31054 37502 31106
rect 36318 31042 36370 31054
rect 32062 30994 32114 31006
rect 28130 30942 28142 30994
rect 28194 30942 28206 30994
rect 32062 30930 32114 30942
rect 32174 30994 32226 31006
rect 32174 30930 32226 30942
rect 32510 30994 32562 31006
rect 32510 30930 32562 30942
rect 33406 30994 33458 31006
rect 33406 30930 33458 30942
rect 35646 30994 35698 31006
rect 36754 30942 36766 30994
rect 36818 30942 36830 30994
rect 41570 30942 41582 30994
rect 41634 30942 41646 30994
rect 35646 30930 35698 30942
rect 33630 30882 33682 30894
rect 30930 30830 30942 30882
rect 30994 30830 31006 30882
rect 39554 30830 39566 30882
rect 39618 30830 39630 30882
rect 42354 30830 42366 30882
rect 42418 30830 42430 30882
rect 44482 30830 44494 30882
rect 44546 30830 44558 30882
rect 33630 30818 33682 30830
rect 35758 30770 35810 30782
rect 35758 30706 35810 30718
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 42030 30434 42082 30446
rect 42030 30370 42082 30382
rect 42366 30434 42418 30446
rect 42366 30370 42418 30382
rect 36094 30322 36146 30334
rect 40350 30322 40402 30334
rect 38546 30270 38558 30322
rect 38610 30270 38622 30322
rect 36094 30258 36146 30270
rect 40350 30258 40402 30270
rect 78206 30322 78258 30334
rect 78206 30258 78258 30270
rect 36206 30210 36258 30222
rect 36206 30146 36258 30158
rect 37774 30210 37826 30222
rect 41022 30210 41074 30222
rect 38434 30158 38446 30210
rect 38498 30158 38510 30210
rect 39890 30158 39902 30210
rect 39954 30158 39966 30210
rect 37774 30146 37826 30158
rect 41022 30146 41074 30158
rect 42254 30210 42306 30222
rect 42254 30146 42306 30158
rect 40462 30098 40514 30110
rect 39778 30046 39790 30098
rect 39842 30046 39854 30098
rect 40462 30034 40514 30046
rect 40686 29986 40738 29998
rect 39554 29934 39566 29986
rect 39618 29934 39630 29986
rect 40686 29922 40738 29934
rect 42366 29986 42418 29998
rect 42366 29922 42418 29934
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 31390 29650 31442 29662
rect 31390 29586 31442 29598
rect 37102 29650 37154 29662
rect 37102 29586 37154 29598
rect 37886 29650 37938 29662
rect 37886 29586 37938 29598
rect 38558 29650 38610 29662
rect 38558 29586 38610 29598
rect 38110 29538 38162 29550
rect 38110 29474 38162 29486
rect 40014 29538 40066 29550
rect 40014 29474 40066 29486
rect 78206 29538 78258 29550
rect 78206 29474 78258 29486
rect 33518 29426 33570 29438
rect 33518 29362 33570 29374
rect 35198 29426 35250 29438
rect 36206 29426 36258 29438
rect 39678 29426 39730 29438
rect 35634 29374 35646 29426
rect 35698 29374 35710 29426
rect 36642 29374 36654 29426
rect 36706 29374 36718 29426
rect 39442 29374 39454 29426
rect 39506 29374 39518 29426
rect 35198 29362 35250 29374
rect 36206 29362 36258 29374
rect 39678 29362 39730 29374
rect 36430 29314 36482 29326
rect 36430 29250 36482 29262
rect 36990 29314 37042 29326
rect 36990 29250 37042 29262
rect 39902 29314 39954 29326
rect 39902 29250 39954 29262
rect 31278 29202 31330 29214
rect 31278 29138 31330 29150
rect 31614 29202 31666 29214
rect 31614 29138 31666 29150
rect 33406 29202 33458 29214
rect 33406 29138 33458 29150
rect 33742 29202 33794 29214
rect 33742 29138 33794 29150
rect 33854 29202 33906 29214
rect 33854 29138 33906 29150
rect 35086 29202 35138 29214
rect 35086 29138 35138 29150
rect 35422 29202 35474 29214
rect 35422 29138 35474 29150
rect 36094 29202 36146 29214
rect 36094 29138 36146 29150
rect 37774 29202 37826 29214
rect 37774 29138 37826 29150
rect 38446 29202 38498 29214
rect 38446 29138 38498 29150
rect 38782 29202 38834 29214
rect 39442 29150 39454 29202
rect 39506 29150 39518 29202
rect 38782 29138 38834 29150
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 36206 28866 36258 28878
rect 36206 28802 36258 28814
rect 38670 28754 38722 28766
rect 30146 28702 30158 28754
rect 30210 28702 30222 28754
rect 32274 28702 32286 28754
rect 32338 28702 32350 28754
rect 33394 28702 33406 28754
rect 33458 28702 33470 28754
rect 35522 28702 35534 28754
rect 35586 28702 35598 28754
rect 35970 28702 35982 28754
rect 36034 28702 36046 28754
rect 37874 28702 37886 28754
rect 37938 28702 37950 28754
rect 39778 28702 39790 28754
rect 39842 28702 39854 28754
rect 41906 28702 41918 28754
rect 41970 28702 41982 28754
rect 38670 28690 38722 28702
rect 29362 28590 29374 28642
rect 29426 28590 29438 28642
rect 32610 28590 32622 28642
rect 32674 28590 32686 28642
rect 35858 28590 35870 28642
rect 35922 28590 35934 28642
rect 38210 28590 38222 28642
rect 38274 28590 38286 28642
rect 39106 28590 39118 28642
rect 39170 28590 39182 28642
rect 78206 28418 78258 28430
rect 78206 28354 78258 28366
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 40910 28082 40962 28094
rect 40910 28018 40962 28030
rect 41022 27970 41074 27982
rect 34738 27918 34750 27970
rect 34802 27918 34814 27970
rect 38210 27918 38222 27970
rect 38274 27918 38286 27970
rect 41022 27906 41074 27918
rect 32274 27806 32286 27858
rect 32338 27806 32350 27858
rect 33954 27806 33966 27858
rect 34018 27806 34030 27858
rect 37538 27806 37550 27858
rect 37602 27806 37614 27858
rect 31502 27746 31554 27758
rect 32162 27694 32174 27746
rect 32226 27694 32238 27746
rect 36866 27694 36878 27746
rect 36930 27694 36942 27746
rect 40338 27694 40350 27746
rect 40402 27694 40414 27746
rect 31502 27682 31554 27694
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 37326 27298 37378 27310
rect 37326 27234 37378 27246
rect 78206 27186 78258 27198
rect 37090 27134 37102 27186
rect 37154 27134 37166 27186
rect 78206 27122 78258 27134
rect 36978 27022 36990 27074
rect 37042 27022 37054 27074
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 78206 20242 78258 20254
rect 78206 20178 78258 20190
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 78206 19346 78258 19358
rect 78206 19282 78258 19294
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 78206 17442 78258 17454
rect 78206 17378 78258 17390
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 78206 16994 78258 17006
rect 78206 16930 78258 16942
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 78206 15874 78258 15886
rect 78206 15810 78258 15822
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 35198 3330 35250 3342
rect 35198 3266 35250 3278
rect 38558 3330 38610 3342
rect 38558 3266 38610 3278
rect 48638 3330 48690 3342
rect 48638 3266 48690 3278
rect 49982 3330 50034 3342
rect 49982 3266 50034 3278
rect 59390 3330 59442 3342
rect 59390 3266 59442 3278
rect 62750 3330 62802 3342
rect 62750 3266 62802 3278
rect 63422 3330 63474 3342
rect 63422 3266 63474 3278
rect 67454 3330 67506 3342
rect 67454 3266 67506 3278
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
<< via1 >>
rect 50430 77198 50482 77250
rect 51214 77198 51266 77250
rect 49758 76974 49810 77026
rect 50318 76974 50370 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 25790 76638 25842 76690
rect 30494 76638 30546 76690
rect 34526 76638 34578 76690
rect 50318 76638 50370 76690
rect 51214 76638 51266 76690
rect 58046 76638 58098 76690
rect 58830 76638 58882 76690
rect 59390 76638 59442 76690
rect 60062 76638 60114 76690
rect 60734 76638 60786 76690
rect 49982 76414 50034 76466
rect 35198 76302 35250 76354
rect 35982 76302 36034 76354
rect 47630 76302 47682 76354
rect 56702 76302 56754 76354
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 50206 75630 50258 75682
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 78206 64542 78258 64594
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 78206 60510 78258 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 78206 59838 78258 59890
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 78206 58158 78258 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 78206 50318 78258 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 47854 49086 47906 49138
rect 44942 48974 44994 49026
rect 45614 48862 45666 48914
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 45614 48414 45666 48466
rect 47630 48414 47682 48466
rect 48750 48414 48802 48466
rect 45838 48302 45890 48354
rect 47742 48302 47794 48354
rect 45950 48190 46002 48242
rect 47406 48190 47458 48242
rect 48190 48190 48242 48242
rect 49086 48190 49138 48242
rect 50878 48190 50930 48242
rect 75630 48190 75682 48242
rect 47518 48078 47570 48130
rect 49534 48078 49586 48130
rect 49982 48078 50034 48130
rect 50542 48078 50594 48130
rect 51550 48078 51602 48130
rect 53678 48078 53730 48130
rect 75406 48078 75458 48130
rect 49422 47966 49474 48018
rect 77982 47966 78034 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 35870 47518 35922 47570
rect 51550 47518 51602 47570
rect 32958 47406 33010 47458
rect 46398 47406 46450 47458
rect 46734 47406 46786 47458
rect 47854 47406 47906 47458
rect 48078 47406 48130 47458
rect 48302 47406 48354 47458
rect 48862 47406 48914 47458
rect 48974 47406 49026 47458
rect 49198 47406 49250 47458
rect 49422 47406 49474 47458
rect 50206 47406 50258 47458
rect 51886 47406 51938 47458
rect 52782 47406 52834 47458
rect 30606 47294 30658 47346
rect 33742 47294 33794 47346
rect 45502 47294 45554 47346
rect 46286 47294 46338 47346
rect 47070 47294 47122 47346
rect 47742 47294 47794 47346
rect 49870 47294 49922 47346
rect 51438 47294 51490 47346
rect 51774 47294 51826 47346
rect 52670 47294 52722 47346
rect 53342 47294 53394 47346
rect 77870 47294 77922 47346
rect 30382 47182 30434 47234
rect 30494 47182 30546 47234
rect 45614 47182 45666 47234
rect 46622 47182 46674 47234
rect 47406 47182 47458 47234
rect 48638 47182 48690 47234
rect 49982 47182 50034 47234
rect 50542 47182 50594 47234
rect 77646 47182 77698 47234
rect 78206 47182 78258 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 34526 46846 34578 46898
rect 34638 46846 34690 46898
rect 46622 46846 46674 46898
rect 50206 46846 50258 46898
rect 51102 46846 51154 46898
rect 29150 46734 29202 46786
rect 46846 46734 46898 46786
rect 48190 46734 48242 46786
rect 48302 46734 48354 46786
rect 49086 46734 49138 46786
rect 49422 46734 49474 46786
rect 49646 46734 49698 46786
rect 50094 46734 50146 46786
rect 50318 46734 50370 46786
rect 78206 46734 78258 46786
rect 28478 46622 28530 46674
rect 31614 46622 31666 46674
rect 31950 46622 32002 46674
rect 32286 46622 32338 46674
rect 33630 46622 33682 46674
rect 38334 46622 38386 46674
rect 42254 46622 42306 46674
rect 46174 46622 46226 46674
rect 46398 46622 46450 46674
rect 47630 46622 47682 46674
rect 47742 46622 47794 46674
rect 47966 46622 48018 46674
rect 48750 46622 48802 46674
rect 50878 46622 50930 46674
rect 31278 46510 31330 46562
rect 31838 46510 31890 46562
rect 33182 46510 33234 46562
rect 34078 46510 34130 46562
rect 34414 46510 34466 46562
rect 35534 46510 35586 46562
rect 37662 46510 37714 46562
rect 43038 46510 43090 46562
rect 45166 46510 45218 46562
rect 46510 46510 46562 46562
rect 49758 46510 49810 46562
rect 48862 46398 48914 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 37550 46062 37602 46114
rect 47182 46062 47234 46114
rect 47518 46062 47570 46114
rect 48414 46062 48466 46114
rect 32062 45950 32114 46002
rect 33070 45950 33122 46002
rect 41134 45950 41186 46002
rect 46846 45950 46898 46002
rect 47630 45950 47682 46002
rect 49422 45950 49474 46002
rect 51102 45950 51154 46002
rect 29262 45838 29314 45890
rect 33294 45838 33346 45890
rect 34414 45838 34466 45890
rect 34638 45838 34690 45890
rect 35086 45838 35138 45890
rect 35646 45838 35698 45890
rect 36990 45838 37042 45890
rect 37214 45838 37266 45890
rect 37438 45838 37490 45890
rect 38334 45838 38386 45890
rect 48302 45838 48354 45890
rect 48638 45838 48690 45890
rect 49086 45838 49138 45890
rect 50206 45838 50258 45890
rect 50654 45838 50706 45890
rect 51998 45838 52050 45890
rect 77646 45838 77698 45890
rect 29934 45726 29986 45778
rect 35534 45726 35586 45778
rect 39006 45726 39058 45778
rect 47966 45726 48018 45778
rect 49310 45726 49362 45778
rect 51438 45726 51490 45778
rect 77422 45726 77474 45778
rect 78206 45726 78258 45778
rect 33630 45614 33682 45666
rect 34078 45614 34130 45666
rect 35422 45614 35474 45666
rect 46958 45614 47010 45666
rect 48078 45614 48130 45666
rect 49870 45614 49922 45666
rect 51550 45614 51602 45666
rect 51662 45614 51714 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 33294 45278 33346 45330
rect 34190 45278 34242 45330
rect 38782 45278 38834 45330
rect 48862 45278 48914 45330
rect 49422 45278 49474 45330
rect 49982 45278 50034 45330
rect 31614 45166 31666 45218
rect 34302 45166 34354 45218
rect 35310 45166 35362 45218
rect 36318 45166 36370 45218
rect 46062 45166 46114 45218
rect 50206 45166 50258 45218
rect 50654 45166 50706 45218
rect 31054 45054 31106 45106
rect 31950 45054 32002 45106
rect 32174 45054 32226 45106
rect 33182 45054 33234 45106
rect 33406 45054 33458 45106
rect 33630 45054 33682 45106
rect 33854 45054 33906 45106
rect 34750 45054 34802 45106
rect 36430 45054 36482 45106
rect 38446 45054 38498 45106
rect 38894 45054 38946 45106
rect 39342 45054 39394 45106
rect 39566 45054 39618 45106
rect 45838 45054 45890 45106
rect 46398 45054 46450 45106
rect 47070 45054 47122 45106
rect 47966 45054 48018 45106
rect 49870 45054 49922 45106
rect 51438 45054 51490 45106
rect 52110 45054 52162 45106
rect 75630 45054 75682 45106
rect 30942 44942 30994 44994
rect 45950 44942 46002 44994
rect 47854 44942 47906 44994
rect 54238 44942 54290 44994
rect 75406 44942 75458 44994
rect 77982 44942 78034 44994
rect 30606 44830 30658 44882
rect 31726 44830 31778 44882
rect 37886 44830 37938 44882
rect 38670 44830 38722 44882
rect 39230 44830 39282 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 35534 44494 35586 44546
rect 46398 44494 46450 44546
rect 49870 44494 49922 44546
rect 50318 44494 50370 44546
rect 51886 44494 51938 44546
rect 39790 44382 39842 44434
rect 44270 44382 44322 44434
rect 44830 44382 44882 44434
rect 51326 44382 51378 44434
rect 53342 44382 53394 44434
rect 34638 44270 34690 44322
rect 34750 44270 34802 44322
rect 35086 44270 35138 44322
rect 39006 44270 39058 44322
rect 39230 44270 39282 44322
rect 39566 44270 39618 44322
rect 39902 44270 39954 44322
rect 41470 44270 41522 44322
rect 45278 44270 45330 44322
rect 45838 44270 45890 44322
rect 46510 44270 46562 44322
rect 50430 44270 50482 44322
rect 51102 44270 51154 44322
rect 51998 44270 52050 44322
rect 34862 44158 34914 44210
rect 38670 44158 38722 44210
rect 42142 44158 42194 44210
rect 45390 44158 45442 44210
rect 45614 44158 45666 44210
rect 49758 44158 49810 44210
rect 51438 44158 51490 44210
rect 52670 44158 52722 44210
rect 52782 44158 52834 44210
rect 39118 44046 39170 44098
rect 44942 44046 44994 44098
rect 46398 44046 46450 44098
rect 50318 44046 50370 44098
rect 51886 44046 51938 44098
rect 53006 44046 53058 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 78206 43710 78258 43762
rect 34302 43598 34354 43650
rect 40238 43598 40290 43650
rect 40350 43598 40402 43650
rect 43374 43598 43426 43650
rect 31054 43486 31106 43538
rect 31278 43486 31330 43538
rect 31726 43486 31778 43538
rect 31950 43486 32002 43538
rect 33966 43486 34018 43538
rect 37886 43486 37938 43538
rect 38446 43486 38498 43538
rect 39342 43486 39394 43538
rect 39790 43486 39842 43538
rect 42590 43486 42642 43538
rect 51326 43486 51378 43538
rect 45502 43374 45554 43426
rect 46286 43374 46338 43426
rect 50878 43374 50930 43426
rect 30718 43262 30770 43314
rect 30830 43262 30882 43314
rect 31614 43262 31666 43314
rect 38110 43262 38162 43314
rect 38558 43262 38610 43314
rect 38670 43262 38722 43314
rect 39566 43262 39618 43314
rect 39902 43262 39954 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 37886 42926 37938 42978
rect 47406 42926 47458 42978
rect 51102 42926 51154 42978
rect 51326 42926 51378 42978
rect 51886 42926 51938 42978
rect 52782 42926 52834 42978
rect 29934 42814 29986 42866
rect 32062 42814 32114 42866
rect 36318 42814 36370 42866
rect 37214 42814 37266 42866
rect 42030 42814 42082 42866
rect 50542 42814 50594 42866
rect 29262 42702 29314 42754
rect 33294 42702 33346 42754
rect 36430 42702 36482 42754
rect 37438 42702 37490 42754
rect 37662 42702 37714 42754
rect 38782 42702 38834 42754
rect 45950 42702 46002 42754
rect 46846 42702 46898 42754
rect 52670 42702 52722 42754
rect 33070 42590 33122 42642
rect 33518 42590 33570 42642
rect 33742 42590 33794 42642
rect 47182 42590 47234 42642
rect 50654 42590 50706 42642
rect 51550 42590 51602 42642
rect 51662 42590 51714 42642
rect 33854 42478 33906 42530
rect 38334 42478 38386 42530
rect 45614 42478 45666 42530
rect 46286 42478 46338 42530
rect 47742 42478 47794 42530
rect 50430 42478 50482 42530
rect 52782 42478 52834 42530
rect 53454 42478 53506 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 31166 42142 31218 42194
rect 44606 42142 44658 42194
rect 49086 42030 49138 42082
rect 51438 42030 51490 42082
rect 28030 41918 28082 41970
rect 31726 41918 31778 41970
rect 32398 41918 32450 41970
rect 38558 41918 38610 41970
rect 38894 41918 38946 41970
rect 39118 41918 39170 41970
rect 39342 41918 39394 41970
rect 39566 41918 39618 41970
rect 40798 41918 40850 41970
rect 41134 41918 41186 41970
rect 41358 41918 41410 41970
rect 44942 41918 44994 41970
rect 45278 41918 45330 41970
rect 48750 41918 48802 41970
rect 50654 41918 50706 41970
rect 75630 41918 75682 41970
rect 28702 41806 28754 41858
rect 30830 41806 30882 41858
rect 32174 41806 32226 41858
rect 33518 41806 33570 41858
rect 41022 41806 41074 41858
rect 46062 41806 46114 41858
rect 48190 41806 48242 41858
rect 53566 41806 53618 41858
rect 75294 41806 75346 41858
rect 77982 41806 78034 41858
rect 31502 41694 31554 41746
rect 32062 41694 32114 41746
rect 39678 41694 39730 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 30606 41358 30658 41410
rect 30942 41358 30994 41410
rect 33406 41358 33458 41410
rect 38334 41358 38386 41410
rect 38558 41358 38610 41410
rect 38670 41358 38722 41410
rect 45614 41358 45666 41410
rect 45950 41358 46002 41410
rect 32398 41246 32450 41298
rect 39118 41246 39170 41298
rect 41246 41246 41298 41298
rect 49310 41246 49362 41298
rect 30718 41134 30770 41186
rect 31166 41134 31218 41186
rect 32958 41134 33010 41186
rect 37438 41134 37490 41186
rect 38110 41134 38162 41186
rect 42030 41134 42082 41186
rect 42814 41134 42866 41186
rect 43486 41134 43538 41186
rect 44158 41134 44210 41186
rect 46398 41134 46450 41186
rect 32510 41022 32562 41074
rect 32734 41022 32786 41074
rect 37662 41022 37714 41074
rect 43038 41022 43090 41074
rect 43822 41022 43874 41074
rect 45838 41022 45890 41074
rect 47182 41022 47234 41074
rect 77646 41022 77698 41074
rect 77870 41022 77922 41074
rect 78206 41022 78258 41074
rect 43934 40910 43986 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 31726 40574 31778 40626
rect 41470 40574 41522 40626
rect 41694 40574 41746 40626
rect 46398 40574 46450 40626
rect 75294 40574 75346 40626
rect 34302 40462 34354 40514
rect 34638 40462 34690 40514
rect 37102 40462 37154 40514
rect 39006 40462 39058 40514
rect 42254 40462 42306 40514
rect 43374 40462 43426 40514
rect 47966 40462 48018 40514
rect 49534 40462 49586 40514
rect 77310 40462 77362 40514
rect 31614 40350 31666 40402
rect 31838 40350 31890 40402
rect 32174 40350 32226 40402
rect 37886 40350 37938 40402
rect 39230 40350 39282 40402
rect 42702 40350 42754 40402
rect 47742 40350 47794 40402
rect 48862 40350 48914 40402
rect 75630 40350 75682 40402
rect 34974 40238 35026 40290
rect 45502 40238 45554 40290
rect 46510 40238 46562 40290
rect 51662 40238 51714 40290
rect 42030 40126 42082 40178
rect 46174 40126 46226 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 30382 39790 30434 39842
rect 30606 39790 30658 39842
rect 31166 39790 31218 39842
rect 31502 39790 31554 39842
rect 32062 39790 32114 39842
rect 32398 39790 32450 39842
rect 32958 39790 33010 39842
rect 43598 39790 43650 39842
rect 33070 39678 33122 39730
rect 39342 39678 39394 39730
rect 42926 39678 42978 39730
rect 30830 39566 30882 39618
rect 31726 39566 31778 39618
rect 32622 39566 32674 39618
rect 35758 39566 35810 39618
rect 42142 39566 42194 39618
rect 43262 39566 43314 39618
rect 30270 39454 30322 39506
rect 33182 39454 33234 39506
rect 41470 39454 41522 39506
rect 35422 39342 35474 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 35086 39006 35138 39058
rect 35422 39006 35474 39058
rect 37774 39006 37826 39058
rect 30382 38894 30434 38946
rect 37102 38894 37154 38946
rect 41134 38894 41186 38946
rect 29710 38782 29762 38834
rect 37998 38782 38050 38834
rect 39454 38782 39506 38834
rect 40350 38782 40402 38834
rect 40910 38782 40962 38834
rect 32510 38670 32562 38722
rect 36990 38670 37042 38722
rect 39790 38670 39842 38722
rect 41246 38670 41298 38722
rect 37326 38558 37378 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 35534 38222 35586 38274
rect 30046 38110 30098 38162
rect 31502 38110 31554 38162
rect 39566 38110 39618 38162
rect 31614 37998 31666 38050
rect 35758 37998 35810 38050
rect 35982 37998 36034 38050
rect 36990 37998 37042 38050
rect 30158 37886 30210 37938
rect 30382 37886 30434 37938
rect 30718 37886 30770 37938
rect 35422 37886 35474 37938
rect 36430 37774 36482 37826
rect 78206 37774 78258 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 38558 37438 38610 37490
rect 40350 37438 40402 37490
rect 29710 37326 29762 37378
rect 29038 37214 29090 37266
rect 34750 37214 34802 37266
rect 37998 37214 38050 37266
rect 39454 37214 39506 37266
rect 39566 37214 39618 37266
rect 39678 37214 39730 37266
rect 40126 37214 40178 37266
rect 31838 37102 31890 37154
rect 35534 37102 35586 37154
rect 37662 37102 37714 37154
rect 38222 36990 38274 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 36990 36654 37042 36706
rect 37998 36654 38050 36706
rect 38110 36654 38162 36706
rect 38334 36654 38386 36706
rect 41022 36654 41074 36706
rect 34302 36542 34354 36594
rect 36430 36542 36482 36594
rect 38894 36542 38946 36594
rect 42814 36542 42866 36594
rect 32510 36430 32562 36482
rect 33630 36430 33682 36482
rect 38446 36430 38498 36482
rect 39118 36430 39170 36482
rect 39678 36430 39730 36482
rect 40014 36430 40066 36482
rect 40350 36430 40402 36482
rect 40686 36430 40738 36482
rect 41134 36430 41186 36482
rect 41358 36430 41410 36482
rect 41582 36430 41634 36482
rect 41806 36430 41858 36482
rect 42590 36430 42642 36482
rect 37102 36318 37154 36370
rect 37326 36318 37378 36370
rect 39342 36318 39394 36370
rect 42926 36318 42978 36370
rect 32174 36206 32226 36258
rect 39902 36206 39954 36258
rect 40238 36206 40290 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 43262 35758 43314 35810
rect 42478 35646 42530 35698
rect 45390 35534 45442 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 42926 35086 42978 35138
rect 32062 34974 32114 35026
rect 41470 34974 41522 35026
rect 42590 34974 42642 35026
rect 29150 34862 29202 34914
rect 38670 34862 38722 34914
rect 42254 34862 42306 34914
rect 29934 34750 29986 34802
rect 32398 34750 32450 34802
rect 39342 34750 39394 34802
rect 32510 34638 32562 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 31390 34302 31442 34354
rect 35422 34302 35474 34354
rect 37102 34302 37154 34354
rect 41246 34302 41298 34354
rect 32398 34190 32450 34242
rect 32510 34190 32562 34242
rect 35086 34190 35138 34242
rect 37438 34190 37490 34242
rect 39790 34190 39842 34242
rect 40910 34190 40962 34242
rect 42702 34190 42754 34242
rect 43262 34190 43314 34242
rect 31502 34078 31554 34130
rect 33406 34078 33458 34130
rect 39902 34078 39954 34130
rect 40238 34078 40290 34130
rect 42142 34078 42194 34130
rect 42366 34078 42418 34130
rect 43038 34078 43090 34130
rect 43150 33966 43202 34018
rect 31390 33854 31442 33906
rect 31726 33854 31778 33906
rect 32398 33854 32450 33906
rect 33630 33854 33682 33906
rect 33854 33854 33906 33906
rect 33966 33854 34018 33906
rect 40126 33854 40178 33906
rect 41806 33854 41858 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 33182 33518 33234 33570
rect 31390 33406 31442 33458
rect 34750 33406 34802 33458
rect 37438 33406 37490 33458
rect 40574 33406 40626 33458
rect 31278 33294 31330 33346
rect 32174 33294 32226 33346
rect 32734 33294 32786 33346
rect 33966 33294 34018 33346
rect 34974 33294 35026 33346
rect 36206 33294 36258 33346
rect 39230 33294 39282 33346
rect 31614 33182 31666 33234
rect 31838 33182 31890 33234
rect 32286 33182 32338 33234
rect 32510 33182 32562 33234
rect 34078 33182 34130 33234
rect 35646 33182 35698 33234
rect 37774 33182 37826 33234
rect 44046 33182 44098 33234
rect 35982 33070 36034 33122
rect 37550 33070 37602 33122
rect 43822 33070 43874 33122
rect 43934 33070 43986 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 34638 32622 34690 32674
rect 30942 32510 30994 32562
rect 31950 32510 32002 32562
rect 32174 32510 32226 32562
rect 38334 32510 38386 32562
rect 39790 32510 39842 32562
rect 44158 32510 44210 32562
rect 31054 32398 31106 32450
rect 40014 32398 40066 32450
rect 41358 32398 41410 32450
rect 43486 32398 43538 32450
rect 30718 32286 30770 32338
rect 32510 32286 32562 32338
rect 40350 32286 40402 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 30718 31950 30770 32002
rect 39678 31950 39730 32002
rect 43150 31950 43202 32002
rect 45054 31950 45106 32002
rect 31502 31838 31554 31890
rect 33630 31838 33682 31890
rect 43486 31838 43538 31890
rect 43598 31838 43650 31890
rect 34414 31726 34466 31778
rect 36990 31726 37042 31778
rect 37998 31726 38050 31778
rect 39118 31726 39170 31778
rect 39566 31726 39618 31778
rect 42142 31726 42194 31778
rect 43262 31726 43314 31778
rect 44830 31726 44882 31778
rect 37102 31614 37154 31666
rect 38558 31614 38610 31666
rect 41022 31614 41074 31666
rect 42030 31614 42082 31666
rect 30494 31502 30546 31554
rect 30606 31502 30658 31554
rect 37214 31502 37266 31554
rect 39006 31502 39058 31554
rect 45390 31502 45442 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 32398 31166 32450 31218
rect 33070 31166 33122 31218
rect 34302 31166 34354 31218
rect 35870 31166 35922 31218
rect 36094 31166 36146 31218
rect 28814 31054 28866 31106
rect 33966 31054 34018 31106
rect 36318 31054 36370 31106
rect 37438 31054 37490 31106
rect 28142 30942 28194 30994
rect 32062 30942 32114 30994
rect 32174 30942 32226 30994
rect 32510 30942 32562 30994
rect 33406 30942 33458 30994
rect 35646 30942 35698 30994
rect 36766 30942 36818 30994
rect 41582 30942 41634 30994
rect 30942 30830 30994 30882
rect 33630 30830 33682 30882
rect 39566 30830 39618 30882
rect 42366 30830 42418 30882
rect 44494 30830 44546 30882
rect 35758 30718 35810 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 42030 30382 42082 30434
rect 42366 30382 42418 30434
rect 36094 30270 36146 30322
rect 38558 30270 38610 30322
rect 40350 30270 40402 30322
rect 78206 30270 78258 30322
rect 36206 30158 36258 30210
rect 37774 30158 37826 30210
rect 38446 30158 38498 30210
rect 39902 30158 39954 30210
rect 41022 30158 41074 30210
rect 42254 30158 42306 30210
rect 39790 30046 39842 30098
rect 40462 30046 40514 30098
rect 39566 29934 39618 29986
rect 40686 29934 40738 29986
rect 42366 29934 42418 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 31390 29598 31442 29650
rect 37102 29598 37154 29650
rect 37886 29598 37938 29650
rect 38558 29598 38610 29650
rect 38110 29486 38162 29538
rect 40014 29486 40066 29538
rect 78206 29486 78258 29538
rect 33518 29374 33570 29426
rect 35198 29374 35250 29426
rect 35646 29374 35698 29426
rect 36206 29374 36258 29426
rect 36654 29374 36706 29426
rect 39454 29374 39506 29426
rect 39678 29374 39730 29426
rect 36430 29262 36482 29314
rect 36990 29262 37042 29314
rect 39902 29262 39954 29314
rect 31278 29150 31330 29202
rect 31614 29150 31666 29202
rect 33406 29150 33458 29202
rect 33742 29150 33794 29202
rect 33854 29150 33906 29202
rect 35086 29150 35138 29202
rect 35422 29150 35474 29202
rect 36094 29150 36146 29202
rect 37774 29150 37826 29202
rect 38446 29150 38498 29202
rect 38782 29150 38834 29202
rect 39454 29150 39506 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 36206 28814 36258 28866
rect 30158 28702 30210 28754
rect 32286 28702 32338 28754
rect 33406 28702 33458 28754
rect 35534 28702 35586 28754
rect 35982 28702 36034 28754
rect 37886 28702 37938 28754
rect 38670 28702 38722 28754
rect 39790 28702 39842 28754
rect 41918 28702 41970 28754
rect 29374 28590 29426 28642
rect 32622 28590 32674 28642
rect 35870 28590 35922 28642
rect 38222 28590 38274 28642
rect 39118 28590 39170 28642
rect 78206 28366 78258 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 40910 28030 40962 28082
rect 34750 27918 34802 27970
rect 38222 27918 38274 27970
rect 41022 27918 41074 27970
rect 32286 27806 32338 27858
rect 33966 27806 34018 27858
rect 37550 27806 37602 27858
rect 31502 27694 31554 27746
rect 32174 27694 32226 27746
rect 36878 27694 36930 27746
rect 40350 27694 40402 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 37326 27246 37378 27298
rect 37102 27134 37154 27186
rect 78206 27134 78258 27186
rect 36990 27022 37042 27074
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 78206 20190 78258 20242
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 78206 19294 78258 19346
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 78206 17390 78258 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 78206 16942 78258 16994
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 78206 15822 78258 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 35198 3278 35250 3330
rect 38558 3278 38610 3330
rect 48638 3278 48690 3330
rect 49982 3278 50034 3330
rect 59390 3278 59442 3330
rect 62750 3278 62802 3330
rect 63422 3278 63474 3330
rect 67454 3278 67506 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 25536 79200 25648 80000
rect 30240 79200 30352 80000
rect 34272 79200 34384 80000
rect 34944 79200 35056 80000
rect 35616 79200 35728 80000
rect 47040 79200 47152 80000
rect 49728 79200 49840 80000
rect 50400 79200 50512 80000
rect 56448 79200 56560 80000
rect 57792 79200 57904 80000
rect 58464 79200 58576 80000
rect 59136 79200 59248 80000
rect 59808 79200 59920 80000
rect 60480 79200 60592 80000
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 25564 76692 25620 79200
rect 25788 76692 25844 76702
rect 25564 76690 25844 76692
rect 25564 76638 25790 76690
rect 25842 76638 25844 76690
rect 25564 76636 25844 76638
rect 30268 76692 30324 79200
rect 30492 76692 30548 76702
rect 30268 76690 30548 76692
rect 30268 76638 30494 76690
rect 30546 76638 30548 76690
rect 30268 76636 30548 76638
rect 34300 76692 34356 79200
rect 34524 76692 34580 76702
rect 34300 76690 34580 76692
rect 34300 76638 34526 76690
rect 34578 76638 34580 76690
rect 34300 76636 34580 76638
rect 25788 76626 25844 76636
rect 30492 76626 30548 76636
rect 34524 76626 34580 76636
rect 34972 76356 35028 79200
rect 35644 77700 35700 79200
rect 35644 77644 36036 77700
rect 35196 76356 35252 76366
rect 34972 76354 35252 76356
rect 34972 76302 35198 76354
rect 35250 76302 35252 76354
rect 34972 76300 35252 76302
rect 35196 76290 35252 76300
rect 35980 76354 36036 77644
rect 35980 76302 35982 76354
rect 36034 76302 36036 76354
rect 35980 76290 36036 76302
rect 47068 76356 47124 79200
rect 49756 77026 49812 79200
rect 50428 77250 50484 79200
rect 50428 77198 50430 77250
rect 50482 77198 50484 77250
rect 50428 77186 50484 77198
rect 51212 77250 51268 77262
rect 51212 77198 51214 77250
rect 51266 77198 51268 77250
rect 49756 76974 49758 77026
rect 49810 76974 49812 77026
rect 49756 76962 49812 76974
rect 50316 77026 50372 77038
rect 50316 76974 50318 77026
rect 50370 76974 50372 77026
rect 50316 76690 50372 76974
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50316 76638 50318 76690
rect 50370 76638 50372 76690
rect 50316 76626 50372 76638
rect 51212 76690 51268 77198
rect 51212 76638 51214 76690
rect 51266 76638 51268 76690
rect 51212 76626 51268 76638
rect 49980 76468 50036 76478
rect 49980 76466 50260 76468
rect 49980 76414 49982 76466
rect 50034 76414 50260 76466
rect 49980 76412 50260 76414
rect 49980 76402 50036 76412
rect 47628 76356 47684 76366
rect 47068 76354 47684 76356
rect 47068 76302 47630 76354
rect 47682 76302 47684 76354
rect 47068 76300 47684 76302
rect 47628 76290 47684 76300
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 50204 75682 50260 76412
rect 56476 76356 56532 79200
rect 57820 76692 57876 79200
rect 58044 76692 58100 76702
rect 57820 76690 58100 76692
rect 57820 76638 58046 76690
rect 58098 76638 58100 76690
rect 57820 76636 58100 76638
rect 58492 76692 58548 79200
rect 58828 76692 58884 76702
rect 58492 76690 58884 76692
rect 58492 76638 58830 76690
rect 58882 76638 58884 76690
rect 58492 76636 58884 76638
rect 59164 76692 59220 79200
rect 59388 76692 59444 76702
rect 59164 76690 59444 76692
rect 59164 76638 59390 76690
rect 59442 76638 59444 76690
rect 59164 76636 59444 76638
rect 59836 76692 59892 79200
rect 60060 76692 60116 76702
rect 59836 76690 60116 76692
rect 59836 76638 60062 76690
rect 60114 76638 60116 76690
rect 59836 76636 60116 76638
rect 60508 76692 60564 79200
rect 60732 76692 60788 76702
rect 60508 76690 60788 76692
rect 60508 76638 60734 76690
rect 60786 76638 60788 76690
rect 60508 76636 60788 76638
rect 58044 76626 58100 76636
rect 58828 76626 58884 76636
rect 59388 76626 59444 76636
rect 60060 76626 60116 76636
rect 60732 76626 60788 76636
rect 56700 76356 56756 76366
rect 56476 76354 56756 76356
rect 56476 76302 56702 76354
rect 56754 76302 56756 76354
rect 56476 76300 56756 76302
rect 56700 76290 56756 76300
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 50204 75630 50206 75682
rect 50258 75630 50260 75682
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 50204 55468 50260 75630
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 78204 64596 78260 64606
rect 78204 64502 78260 64540
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 78204 60564 78260 60574
rect 78204 60470 78260 60508
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 78204 59892 78260 59902
rect 78204 59798 78260 59836
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 78204 58210 78260 58222
rect 78204 58158 78206 58210
rect 78258 58158 78260 58210
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 78204 57876 78260 58158
rect 78204 57810 78260 57820
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 49532 55412 50260 55468
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 47852 49140 47908 49150
rect 44940 49028 44996 49038
rect 44940 49026 45108 49028
rect 44940 48974 44942 49026
rect 44994 48974 45108 49026
rect 44940 48972 45108 48974
rect 44940 48962 44996 48972
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35868 47570 35924 47582
rect 35868 47518 35870 47570
rect 35922 47518 35924 47570
rect 32956 47458 33012 47470
rect 32956 47406 32958 47458
rect 33010 47406 33012 47458
rect 30604 47346 30660 47358
rect 30604 47294 30606 47346
rect 30658 47294 30660 47346
rect 29148 47236 29204 47246
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 29148 46786 29204 47180
rect 30380 47234 30436 47246
rect 30380 47182 30382 47234
rect 30434 47182 30436 47234
rect 30380 47124 30436 47182
rect 30492 47236 30548 47246
rect 30492 47142 30548 47180
rect 30380 47058 30436 47068
rect 29148 46734 29150 46786
rect 29202 46734 29204 46786
rect 29148 46722 29204 46734
rect 28476 46674 28532 46686
rect 28476 46622 28478 46674
rect 28530 46622 28532 46674
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 28476 45892 28532 46622
rect 28476 45826 28532 45836
rect 29260 45892 29316 45902
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 29260 42754 29316 45836
rect 29932 45778 29988 45790
rect 29932 45726 29934 45778
rect 29986 45726 29988 45778
rect 29932 45332 29988 45726
rect 29932 45266 29988 45276
rect 30604 44882 30660 47294
rect 30940 46732 31668 46788
rect 30940 44994 30996 46732
rect 31612 46674 31668 46732
rect 31612 46622 31614 46674
rect 31666 46622 31668 46674
rect 31612 46610 31668 46622
rect 31948 46674 32004 46686
rect 31948 46622 31950 46674
rect 32002 46622 32004 46674
rect 31276 46564 31332 46574
rect 31052 45108 31108 45118
rect 31276 45108 31332 46508
rect 31836 46562 31892 46574
rect 31836 46510 31838 46562
rect 31890 46510 31892 46562
rect 31612 45332 31668 45342
rect 31612 45218 31668 45276
rect 31612 45166 31614 45218
rect 31666 45166 31668 45218
rect 31612 45154 31668 45166
rect 31052 45106 31332 45108
rect 31052 45054 31054 45106
rect 31106 45054 31332 45106
rect 31052 45052 31332 45054
rect 31836 45108 31892 46510
rect 31948 46564 32004 46622
rect 31948 46498 32004 46508
rect 32284 46674 32340 46686
rect 32284 46622 32286 46674
rect 32338 46622 32340 46674
rect 32060 46002 32116 46014
rect 32060 45950 32062 46002
rect 32114 45950 32116 46002
rect 32060 45892 32116 45950
rect 32284 45892 32340 46622
rect 32396 45892 32452 45902
rect 32060 45836 32396 45892
rect 32396 45826 32452 45836
rect 32172 45668 32228 45678
rect 31948 45108 32004 45118
rect 31836 45106 32004 45108
rect 31836 45054 31950 45106
rect 32002 45054 32004 45106
rect 31836 45052 32004 45054
rect 31052 45042 31108 45052
rect 31948 45042 32004 45052
rect 32172 45106 32228 45612
rect 32172 45054 32174 45106
rect 32226 45054 32228 45106
rect 32172 45042 32228 45054
rect 30940 44942 30942 44994
rect 30994 44942 30996 44994
rect 30604 44830 30606 44882
rect 30658 44830 30660 44882
rect 30604 44818 30660 44830
rect 30828 44884 30884 44894
rect 29932 43316 29988 43326
rect 29932 42866 29988 43260
rect 30716 43316 30772 43326
rect 30716 43222 30772 43260
rect 30828 43314 30884 44828
rect 30940 43652 30996 44942
rect 31724 44884 31780 44894
rect 31724 44790 31780 44828
rect 30940 43540 30996 43596
rect 31052 43540 31108 43550
rect 30940 43538 31108 43540
rect 30940 43486 31054 43538
rect 31106 43486 31108 43538
rect 30940 43484 31108 43486
rect 31052 43474 31108 43484
rect 31276 43540 31332 43550
rect 31724 43540 31780 43550
rect 31276 43538 31780 43540
rect 31276 43486 31278 43538
rect 31330 43486 31726 43538
rect 31778 43486 31780 43538
rect 31276 43484 31780 43486
rect 31276 43474 31332 43484
rect 31724 43474 31780 43484
rect 31948 43540 32004 43550
rect 31948 43538 32116 43540
rect 31948 43486 31950 43538
rect 32002 43486 32116 43538
rect 31948 43484 32116 43486
rect 31948 43474 32004 43484
rect 31612 43316 31668 43326
rect 30828 43262 30830 43314
rect 30882 43262 30884 43314
rect 29932 42814 29934 42866
rect 29986 42814 29988 42866
rect 29932 42802 29988 42814
rect 29260 42702 29262 42754
rect 29314 42702 29316 42754
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 28028 41970 28084 41982
rect 28028 41918 28030 41970
rect 28082 41918 28084 41970
rect 28028 41860 28084 41918
rect 28028 41794 28084 41804
rect 28700 41858 28756 41870
rect 28700 41806 28702 41858
rect 28754 41806 28756 41858
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 28700 41412 28756 41806
rect 29260 41860 29316 42702
rect 30828 42196 30884 43262
rect 31164 43314 31668 43316
rect 31164 43262 31614 43314
rect 31666 43262 31668 43314
rect 31164 43260 31668 43262
rect 31164 42196 31220 43260
rect 31612 43250 31668 43260
rect 32060 42866 32116 43484
rect 32060 42814 32062 42866
rect 32114 42814 32116 42866
rect 32060 42756 32116 42814
rect 32060 42690 32116 42700
rect 32508 42756 32564 42766
rect 30716 42140 30884 42196
rect 30940 42194 31220 42196
rect 30940 42142 31166 42194
rect 31218 42142 31220 42194
rect 30940 42140 31220 42142
rect 29260 41794 29316 41804
rect 29708 41860 29764 41870
rect 28700 41346 28756 41356
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 29708 38834 29764 41804
rect 30604 41412 30660 41422
rect 30604 41318 30660 41356
rect 30716 41186 30772 42140
rect 30828 41972 30884 41982
rect 30828 41858 30884 41916
rect 30828 41806 30830 41858
rect 30882 41806 30884 41858
rect 30828 41794 30884 41806
rect 30940 41410 30996 42140
rect 31164 42130 31220 42140
rect 31724 41972 31780 41982
rect 31724 41878 31780 41916
rect 32396 41972 32452 41982
rect 32172 41858 32228 41870
rect 32172 41806 32174 41858
rect 32226 41806 32228 41858
rect 31500 41748 31556 41758
rect 31500 41654 31556 41692
rect 32060 41748 32116 41758
rect 30940 41358 30942 41410
rect 30994 41358 30996 41410
rect 30940 41346 30996 41358
rect 31164 41412 31220 41422
rect 30716 41134 30718 41186
rect 30770 41134 30772 41186
rect 30380 40292 30436 40302
rect 30380 39842 30436 40236
rect 30716 40292 30772 41134
rect 31164 41186 31220 41356
rect 31164 41134 31166 41186
rect 31218 41134 31220 41186
rect 31164 41122 31220 41134
rect 31724 40628 31780 40638
rect 30716 40226 30772 40236
rect 31052 40626 31780 40628
rect 31052 40574 31726 40626
rect 31778 40574 31780 40626
rect 31052 40572 31780 40574
rect 31052 39956 31108 40572
rect 31724 40562 31780 40572
rect 30380 39790 30382 39842
rect 30434 39790 30436 39842
rect 30380 39778 30436 39790
rect 30604 39900 31108 39956
rect 31164 40404 31220 40414
rect 30604 39842 30660 39900
rect 31164 39844 31220 40348
rect 31612 40402 31668 40414
rect 31612 40350 31614 40402
rect 31666 40350 31668 40402
rect 30604 39790 30606 39842
rect 30658 39790 30660 39842
rect 30604 39778 30660 39790
rect 30828 39842 31220 39844
rect 30828 39790 31166 39842
rect 31218 39790 31220 39842
rect 30828 39788 31220 39790
rect 30828 39618 30884 39788
rect 31164 39778 31220 39788
rect 31500 40068 31556 40078
rect 31500 39842 31556 40012
rect 31500 39790 31502 39842
rect 31554 39790 31556 39842
rect 31500 39778 31556 39790
rect 30828 39566 30830 39618
rect 30882 39566 30884 39618
rect 30828 39554 30884 39566
rect 31612 39620 31668 40350
rect 31836 40402 31892 40414
rect 31836 40350 31838 40402
rect 31890 40350 31892 40402
rect 31724 39620 31780 39630
rect 31612 39618 31780 39620
rect 31612 39566 31726 39618
rect 31778 39566 31780 39618
rect 31612 39564 31780 39566
rect 30268 39506 30324 39518
rect 30268 39454 30270 39506
rect 30322 39454 30324 39506
rect 30268 38948 30324 39454
rect 30380 38948 30436 38958
rect 30268 38946 30436 38948
rect 30268 38894 30382 38946
rect 30434 38894 30436 38946
rect 30268 38892 30436 38894
rect 30380 38882 30436 38892
rect 29708 38782 29710 38834
rect 29762 38782 29764 38834
rect 29708 38770 29764 38782
rect 31724 38668 31780 39564
rect 31500 38612 31780 38668
rect 31836 39508 31892 40350
rect 32060 40404 32116 41692
rect 32172 41412 32228 41806
rect 32172 41346 32228 41356
rect 32396 41298 32452 41916
rect 32396 41246 32398 41298
rect 32450 41246 32452 41298
rect 32396 41234 32452 41246
rect 32508 41074 32564 42700
rect 32956 41860 33012 47406
rect 33740 47348 33796 47358
rect 33740 47346 34580 47348
rect 33740 47294 33742 47346
rect 33794 47294 34580 47346
rect 33740 47292 34580 47294
rect 33740 47282 33796 47292
rect 34524 46898 34580 47292
rect 34524 46846 34526 46898
rect 34578 46846 34580 46898
rect 34524 46834 34580 46846
rect 34636 47124 34692 47134
rect 34636 46898 34692 47068
rect 34636 46846 34638 46898
rect 34690 46846 34692 46898
rect 33628 46676 33684 46686
rect 33628 46674 33796 46676
rect 33628 46622 33630 46674
rect 33682 46622 33796 46674
rect 33628 46620 33796 46622
rect 33628 46610 33684 46620
rect 33068 46564 33124 46574
rect 33068 46002 33124 46508
rect 33068 45950 33070 46002
rect 33122 45950 33124 46002
rect 33068 45108 33124 45950
rect 33180 46562 33236 46574
rect 33180 46510 33182 46562
rect 33234 46510 33236 46562
rect 33180 45668 33236 46510
rect 33292 45892 33348 45902
rect 33348 45836 33460 45892
rect 33292 45798 33348 45836
rect 33180 45602 33236 45612
rect 33292 45330 33348 45342
rect 33292 45278 33294 45330
rect 33346 45278 33348 45330
rect 33180 45108 33236 45118
rect 33068 45106 33236 45108
rect 33068 45054 33182 45106
rect 33234 45054 33236 45106
rect 33068 45052 33236 45054
rect 33180 45042 33236 45052
rect 33292 42754 33348 45278
rect 33404 45106 33460 45836
rect 33628 45666 33684 45678
rect 33628 45614 33630 45666
rect 33682 45614 33684 45666
rect 33628 45332 33684 45614
rect 33628 45266 33684 45276
rect 33740 45332 33796 46620
rect 34076 46564 34132 46574
rect 34412 46564 34468 46574
rect 34076 46562 34468 46564
rect 34076 46510 34078 46562
rect 34130 46510 34414 46562
rect 34466 46510 34468 46562
rect 34076 46508 34468 46510
rect 34076 46498 34132 46508
rect 34412 46498 34468 46508
rect 34636 46116 34692 46846
rect 35532 46564 35588 46574
rect 35532 46562 35700 46564
rect 35532 46510 35534 46562
rect 35586 46510 35700 46562
rect 35532 46508 35700 46510
rect 35532 46498 35588 46508
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34524 46060 34692 46116
rect 34412 45890 34468 45902
rect 34412 45838 34414 45890
rect 34466 45838 34468 45890
rect 34076 45668 34132 45678
rect 34076 45574 34132 45612
rect 34188 45332 34244 45342
rect 33740 45330 34244 45332
rect 33740 45278 34190 45330
rect 34242 45278 34244 45330
rect 33740 45276 34244 45278
rect 33404 45054 33406 45106
rect 33458 45054 33460 45106
rect 33404 45042 33460 45054
rect 33628 45108 33684 45118
rect 33740 45108 33796 45276
rect 34188 45266 34244 45276
rect 34412 45332 34468 45838
rect 34412 45266 34468 45276
rect 34300 45220 34356 45230
rect 34300 45126 34356 45164
rect 33628 45106 33796 45108
rect 33628 45054 33630 45106
rect 33682 45054 33796 45106
rect 33628 45052 33796 45054
rect 33852 45106 33908 45118
rect 33852 45054 33854 45106
rect 33906 45054 33908 45106
rect 33628 45042 33684 45052
rect 33852 44884 33908 45054
rect 33852 44818 33908 44828
rect 33964 45108 34020 45118
rect 33964 43538 34020 45052
rect 34300 43652 34356 43662
rect 34300 43558 34356 43596
rect 33964 43486 33966 43538
rect 34018 43486 34020 43538
rect 33964 43428 34020 43486
rect 33628 43372 34020 43428
rect 33292 42702 33294 42754
rect 33346 42702 33348 42754
rect 33292 42690 33348 42702
rect 33404 42756 33460 42766
rect 32956 41794 33012 41804
rect 33068 42642 33124 42654
rect 33068 42590 33070 42642
rect 33122 42590 33124 42642
rect 32956 41186 33012 41198
rect 32956 41134 32958 41186
rect 33010 41134 33012 41186
rect 32508 41022 32510 41074
rect 32562 41022 32564 41074
rect 32508 41010 32564 41022
rect 32732 41074 32788 41086
rect 32732 41022 32734 41074
rect 32786 41022 32788 41074
rect 32060 40338 32116 40348
rect 32172 40404 32228 40414
rect 32172 40402 32452 40404
rect 32172 40350 32174 40402
rect 32226 40350 32452 40402
rect 32172 40348 32452 40350
rect 32172 40338 32228 40348
rect 32060 40068 32116 40078
rect 32060 39842 32116 40012
rect 32060 39790 32062 39842
rect 32114 39790 32116 39842
rect 32060 39778 32116 39790
rect 32396 39844 32452 40348
rect 32396 39778 32452 39788
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 30044 38164 30100 38174
rect 29708 38162 30100 38164
rect 29708 38110 30046 38162
rect 30098 38110 30100 38162
rect 29708 38108 30100 38110
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 29708 37378 29764 38108
rect 30044 38098 30100 38108
rect 31500 38162 31556 38612
rect 31500 38110 31502 38162
rect 31554 38110 31556 38162
rect 30156 38052 30212 38062
rect 30156 37938 30212 37996
rect 30156 37886 30158 37938
rect 30210 37886 30212 37938
rect 30156 37874 30212 37886
rect 30380 37940 30436 37950
rect 30716 37940 30772 37950
rect 30380 37938 30772 37940
rect 30380 37886 30382 37938
rect 30434 37886 30718 37938
rect 30770 37886 30772 37938
rect 30380 37884 30772 37886
rect 30380 37874 30436 37884
rect 30716 37874 30772 37884
rect 29708 37326 29710 37378
rect 29762 37326 29764 37378
rect 29708 37314 29764 37326
rect 29036 37268 29092 37278
rect 29036 37266 29204 37268
rect 29036 37214 29038 37266
rect 29090 37214 29204 37266
rect 29036 37212 29204 37214
rect 29036 37202 29092 37212
rect 29148 37044 29204 37212
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 29148 34914 29204 36988
rect 29148 34862 29150 34914
rect 29202 34862 29204 34914
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 28140 31892 28196 31902
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 28140 30994 28196 31836
rect 29148 31892 29204 34862
rect 31500 36260 31556 38110
rect 31612 38052 31668 38062
rect 31836 38052 31892 39452
rect 32508 39732 32564 39742
rect 32508 38722 32564 39676
rect 32620 39618 32676 39630
rect 32620 39566 32622 39618
rect 32674 39566 32676 39618
rect 32620 39508 32676 39566
rect 32620 39442 32676 39452
rect 32508 38670 32510 38722
rect 32562 38670 32564 38722
rect 32508 38658 32564 38670
rect 31612 38050 31892 38052
rect 31612 37998 31614 38050
rect 31666 37998 31892 38050
rect 31612 37996 31892 37998
rect 31612 37986 31668 37996
rect 31836 37154 31892 37996
rect 31836 37102 31838 37154
rect 31890 37102 31892 37154
rect 31836 37090 31892 37102
rect 32508 36484 32564 36494
rect 32732 36484 32788 41022
rect 32956 40068 33012 41134
rect 32956 40002 33012 40012
rect 32956 39844 33012 39854
rect 32956 39750 33012 39788
rect 33068 39730 33124 42590
rect 33404 42644 33460 42700
rect 33516 42644 33572 42654
rect 33404 42642 33572 42644
rect 33404 42590 33518 42642
rect 33570 42590 33572 42642
rect 33404 42588 33572 42590
rect 33516 42578 33572 42588
rect 33628 42420 33684 43372
rect 34524 42980 34580 46060
rect 34636 45892 34692 45902
rect 34636 45890 34804 45892
rect 34636 45838 34638 45890
rect 34690 45838 34804 45890
rect 34636 45836 34804 45838
rect 34636 45826 34692 45836
rect 34636 45220 34692 45230
rect 34636 44322 34692 45164
rect 34748 45108 34804 45836
rect 35084 45890 35140 45902
rect 35084 45838 35086 45890
rect 35138 45838 35140 45890
rect 35084 45668 35140 45838
rect 35084 45602 35140 45612
rect 35420 45892 35476 45902
rect 35420 45666 35476 45836
rect 35644 45890 35700 46508
rect 35644 45838 35646 45890
rect 35698 45838 35700 45890
rect 35420 45614 35422 45666
rect 35474 45614 35476 45666
rect 35420 45602 35476 45614
rect 35532 45778 35588 45790
rect 35532 45726 35534 45778
rect 35586 45726 35588 45778
rect 35308 45332 35364 45342
rect 35308 45220 35364 45276
rect 35084 45218 35364 45220
rect 35084 45166 35310 45218
rect 35362 45166 35364 45218
rect 35084 45164 35364 45166
rect 34972 45108 35028 45118
rect 34748 45014 34804 45052
rect 34860 45052 34972 45108
rect 34636 44270 34638 44322
rect 34690 44270 34692 44322
rect 34636 44258 34692 44270
rect 34748 44884 34804 44894
rect 34860 44884 34916 45052
rect 34972 45042 35028 45052
rect 34804 44828 34916 44884
rect 34748 44322 34804 44828
rect 34748 44270 34750 44322
rect 34802 44270 34804 44322
rect 34748 44258 34804 44270
rect 35084 44322 35140 45164
rect 35308 45154 35364 45164
rect 35532 45220 35588 45726
rect 35644 45780 35700 45838
rect 35644 45714 35700 45724
rect 35532 45154 35588 45164
rect 35868 45220 35924 47518
rect 38332 46676 38388 46686
rect 38556 46676 38612 46686
rect 38332 46674 38556 46676
rect 38332 46622 38334 46674
rect 38386 46622 38556 46674
rect 38332 46620 38556 46622
rect 37660 46562 37716 46574
rect 37660 46510 37662 46562
rect 37714 46510 37716 46562
rect 37548 46116 37604 46126
rect 37660 46116 37716 46510
rect 37548 46114 37716 46116
rect 37548 46062 37550 46114
rect 37602 46062 37716 46114
rect 37548 46060 37716 46062
rect 37548 46050 37604 46060
rect 36988 45892 37044 45902
rect 36988 45798 37044 45836
rect 37212 45890 37268 45902
rect 37212 45838 37214 45890
rect 37266 45838 37268 45890
rect 36428 45780 36484 45790
rect 35868 45154 35924 45164
rect 36316 45220 36372 45230
rect 36316 45126 36372 45164
rect 36428 45108 36484 45724
rect 36428 45014 36484 45052
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35532 44548 35588 44558
rect 35532 44454 35588 44492
rect 37212 44548 37268 45838
rect 37436 45892 37492 45902
rect 37436 45890 38276 45892
rect 37436 45838 37438 45890
rect 37490 45838 38276 45890
rect 37436 45836 38276 45838
rect 37436 45826 37492 45836
rect 37212 44482 37268 44492
rect 35084 44270 35086 44322
rect 35138 44270 35140 44322
rect 35084 44258 35140 44270
rect 34860 44210 34916 44222
rect 34860 44158 34862 44210
rect 34914 44158 34916 44210
rect 34860 43652 34916 44158
rect 34860 43586 34916 43596
rect 36316 43540 36372 43550
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34524 42924 35140 42980
rect 33404 42364 33684 42420
rect 33740 42642 33796 42654
rect 33740 42590 33742 42642
rect 33794 42590 33796 42642
rect 33404 41410 33460 42364
rect 33740 41972 33796 42590
rect 33852 42532 33908 42542
rect 33852 42438 33908 42476
rect 33740 41906 33796 41916
rect 34972 42084 35028 42094
rect 33516 41860 33572 41870
rect 33516 41766 33572 41804
rect 33404 41358 33406 41410
rect 33458 41358 33460 41410
rect 33404 41346 33460 41358
rect 34300 40514 34356 40526
rect 34300 40462 34302 40514
rect 34354 40462 34356 40514
rect 34300 40292 34356 40462
rect 34636 40516 34692 40526
rect 34636 40422 34692 40460
rect 34300 40226 34356 40236
rect 34972 40290 35028 42028
rect 34972 40238 34974 40290
rect 35026 40238 35028 40290
rect 34972 40226 35028 40238
rect 33068 39678 33070 39730
rect 33122 39678 33124 39730
rect 33068 39666 33124 39678
rect 33180 39508 33236 39518
rect 33180 39414 33236 39452
rect 35084 39058 35140 42924
rect 36316 42866 36372 43484
rect 36316 42814 36318 42866
rect 36370 42814 36372 42866
rect 36316 42802 36372 42814
rect 37212 42868 37268 42878
rect 37212 42774 37268 42812
rect 36428 42756 36484 42766
rect 36428 42662 36484 42700
rect 37436 42756 37492 42766
rect 37436 42662 37492 42700
rect 37660 42754 37716 42766
rect 37660 42702 37662 42754
rect 37714 42702 37716 42754
rect 37660 42084 37716 42702
rect 37660 42018 37716 42028
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 37436 41186 37492 41198
rect 37436 41134 37438 41186
rect 37490 41134 37492 41186
rect 35756 41076 35812 41086
rect 35756 40516 35812 41020
rect 37436 41076 37492 41134
rect 37436 41010 37492 41020
rect 37660 41076 37716 41086
rect 37772 41076 37828 45836
rect 38220 45220 38276 45836
rect 38332 45890 38388 46620
rect 38556 46610 38612 46620
rect 42028 46676 42084 46686
rect 42252 46676 42308 46686
rect 42084 46674 42308 46676
rect 42084 46622 42254 46674
rect 42306 46622 42308 46674
rect 42084 46620 42308 46622
rect 38332 45838 38334 45890
rect 38386 45838 38388 45890
rect 38332 45826 38388 45838
rect 41132 46002 41188 46014
rect 41132 45950 41134 46002
rect 41186 45950 41188 46002
rect 39004 45780 39060 45790
rect 38780 45778 39060 45780
rect 38780 45726 39006 45778
rect 39058 45726 39060 45778
rect 38780 45724 39060 45726
rect 38780 45330 38836 45724
rect 39004 45714 39060 45724
rect 38780 45278 38782 45330
rect 38834 45278 38836 45330
rect 38780 45266 38836 45278
rect 39564 45332 39620 45342
rect 38220 45164 38500 45220
rect 38444 45106 38500 45164
rect 38444 45054 38446 45106
rect 38498 45054 38500 45106
rect 37884 44882 37940 44894
rect 37884 44830 37886 44882
rect 37938 44830 37940 44882
rect 37884 44324 37940 44830
rect 37884 43538 37940 44268
rect 38444 43876 38500 45054
rect 38892 45108 38948 45118
rect 39340 45108 39396 45118
rect 38892 45106 39396 45108
rect 38892 45054 38894 45106
rect 38946 45054 39342 45106
rect 39394 45054 39396 45106
rect 38892 45052 39396 45054
rect 38892 45042 38948 45052
rect 39340 45042 39396 45052
rect 39564 45106 39620 45276
rect 39564 45054 39566 45106
rect 39618 45054 39620 45106
rect 38668 44884 38724 44894
rect 38668 44790 38724 44828
rect 39228 44882 39284 44894
rect 39228 44830 39230 44882
rect 39282 44830 39284 44882
rect 39004 44660 39060 44670
rect 39004 44322 39060 44604
rect 39004 44270 39006 44322
rect 39058 44270 39060 44322
rect 39004 44258 39060 44270
rect 39228 44548 39284 44830
rect 39564 44660 39620 45054
rect 40348 45332 40404 45342
rect 39564 44594 39620 44604
rect 39788 44884 39844 44894
rect 39228 44322 39284 44492
rect 39788 44434 39844 44828
rect 39788 44382 39790 44434
rect 39842 44382 39844 44434
rect 39788 44370 39844 44382
rect 39228 44270 39230 44322
rect 39282 44270 39284 44322
rect 39228 44258 39284 44270
rect 39564 44324 39620 44334
rect 39564 44230 39620 44268
rect 39900 44322 39956 44334
rect 39900 44270 39902 44322
rect 39954 44270 39956 44322
rect 38444 43810 38500 43820
rect 38668 44210 38724 44222
rect 38668 44158 38670 44210
rect 38722 44158 38724 44210
rect 37884 43486 37886 43538
rect 37938 43486 37940 43538
rect 37884 42980 37940 43486
rect 38444 43652 38500 43662
rect 38444 43538 38500 43596
rect 38444 43486 38446 43538
rect 38498 43486 38500 43538
rect 38444 43428 38500 43486
rect 38668 43540 38724 44158
rect 39116 44098 39172 44110
rect 39116 44046 39118 44098
rect 39170 44046 39172 44098
rect 39116 43652 39172 44046
rect 39452 43652 39508 43662
rect 39900 43652 39956 44270
rect 40236 43652 40292 43662
rect 39116 43596 39396 43652
rect 38724 43484 39284 43540
rect 38668 43474 38724 43484
rect 38220 43372 38500 43428
rect 38108 43314 38164 43326
rect 38108 43262 38110 43314
rect 38162 43262 38164 43314
rect 37884 42978 38052 42980
rect 37884 42926 37886 42978
rect 37938 42926 38052 42978
rect 37884 42924 38052 42926
rect 37884 42914 37940 42924
rect 37996 41188 38052 42924
rect 38108 42756 38164 43262
rect 38108 41412 38164 42700
rect 38220 42868 38276 43372
rect 38556 43316 38612 43326
rect 38220 41636 38276 42812
rect 38444 43314 38612 43316
rect 38444 43262 38558 43314
rect 38610 43262 38612 43314
rect 38444 43260 38612 43262
rect 38332 42530 38388 42542
rect 38332 42478 38334 42530
rect 38386 42478 38388 42530
rect 38332 41972 38388 42478
rect 38332 41906 38388 41916
rect 38444 41860 38500 43260
rect 38556 43250 38612 43260
rect 38668 43314 38724 43326
rect 38668 43262 38670 43314
rect 38722 43262 38724 43314
rect 38668 42980 38724 43262
rect 38556 42924 38724 42980
rect 38556 42196 38612 42924
rect 38556 42130 38612 42140
rect 38780 42754 38836 42766
rect 38780 42702 38782 42754
rect 38834 42702 38836 42754
rect 38556 41972 38612 41982
rect 38780 41972 38836 42702
rect 38556 41970 38836 41972
rect 38556 41918 38558 41970
rect 38610 41918 38836 41970
rect 38556 41916 38836 41918
rect 38556 41906 38612 41916
rect 38444 41794 38500 41804
rect 38220 41580 38500 41636
rect 38332 41412 38388 41422
rect 38108 41410 38388 41412
rect 38108 41358 38334 41410
rect 38386 41358 38388 41410
rect 38108 41356 38388 41358
rect 38444 41412 38500 41580
rect 38556 41412 38612 41422
rect 38444 41410 38612 41412
rect 38444 41358 38558 41410
rect 38610 41358 38612 41410
rect 38444 41356 38612 41358
rect 38332 41346 38388 41356
rect 38556 41346 38612 41356
rect 38668 41412 38724 41422
rect 38668 41318 38724 41356
rect 38108 41188 38164 41198
rect 37996 41186 38164 41188
rect 37996 41134 38110 41186
rect 38162 41134 38164 41186
rect 37996 41132 38164 41134
rect 38108 41122 38164 41132
rect 38780 41188 38836 41916
rect 38892 42532 38948 42542
rect 38892 41970 38948 42476
rect 38892 41918 38894 41970
rect 38946 41918 38948 41970
rect 38892 41906 38948 41918
rect 39116 42084 39172 42094
rect 39116 41970 39172 42028
rect 39116 41918 39118 41970
rect 39170 41918 39172 41970
rect 39116 41906 39172 41918
rect 39228 41972 39284 43484
rect 39340 43538 39396 43596
rect 39508 43596 39844 43652
rect 39452 43586 39508 43596
rect 39340 43486 39342 43538
rect 39394 43486 39396 43538
rect 39340 43474 39396 43486
rect 39788 43538 39844 43596
rect 39788 43486 39790 43538
rect 39842 43486 39844 43538
rect 39788 43474 39844 43486
rect 39900 43650 40292 43652
rect 39900 43598 40238 43650
rect 40290 43598 40292 43650
rect 39900 43596 40292 43598
rect 39900 43540 39956 43596
rect 40236 43586 40292 43596
rect 40348 43650 40404 45276
rect 41132 45332 41188 45950
rect 41132 45266 41188 45276
rect 41468 44324 41524 44334
rect 42028 44324 42084 46620
rect 42252 46610 42308 46620
rect 43036 46564 43092 46574
rect 43036 46470 43092 46508
rect 41468 44322 42084 44324
rect 41468 44270 41470 44322
rect 41522 44270 42084 44322
rect 41468 44268 42084 44270
rect 41468 44258 41524 44268
rect 40348 43598 40350 43650
rect 40402 43598 40404 43650
rect 39900 43474 39956 43484
rect 39564 43316 39620 43326
rect 39452 43314 39620 43316
rect 39452 43262 39566 43314
rect 39618 43262 39620 43314
rect 39452 43260 39620 43262
rect 39340 41972 39396 41982
rect 39228 41970 39396 41972
rect 39228 41918 39342 41970
rect 39394 41918 39396 41970
rect 39228 41916 39396 41918
rect 39116 41300 39172 41310
rect 39228 41300 39284 41916
rect 39340 41906 39396 41916
rect 39452 41412 39508 43260
rect 39564 43250 39620 43260
rect 39900 43314 39956 43326
rect 39900 43262 39902 43314
rect 39954 43262 39956 43314
rect 39564 43092 39620 43102
rect 39564 41970 39620 43036
rect 39564 41918 39566 41970
rect 39618 41918 39620 41970
rect 39564 41906 39620 41918
rect 39452 41346 39508 41356
rect 39676 41746 39732 41758
rect 39676 41694 39678 41746
rect 39730 41694 39732 41746
rect 39116 41298 39284 41300
rect 39116 41246 39118 41298
rect 39170 41246 39284 41298
rect 39116 41244 39284 41246
rect 39116 41234 39172 41244
rect 38780 41122 38836 41132
rect 39564 41188 39620 41198
rect 37660 41074 37828 41076
rect 37660 41022 37662 41074
rect 37714 41022 37828 41074
rect 37660 41020 37828 41022
rect 37660 41010 37716 41020
rect 37772 40628 37828 41020
rect 37772 40562 37828 40572
rect 39228 40628 39284 40638
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35756 39618 35812 40460
rect 37100 40516 37156 40526
rect 37100 40422 37156 40460
rect 39004 40514 39060 40526
rect 39004 40462 39006 40514
rect 39058 40462 39060 40514
rect 37884 40404 37940 40414
rect 37884 40310 37940 40348
rect 39004 40068 39060 40462
rect 39228 40402 39284 40572
rect 39228 40350 39230 40402
rect 39282 40350 39284 40402
rect 39228 40338 39284 40350
rect 39004 40002 39060 40012
rect 35756 39566 35758 39618
rect 35810 39566 35812 39618
rect 35756 39554 35812 39566
rect 39340 39730 39396 39742
rect 39340 39678 39342 39730
rect 39394 39678 39396 39730
rect 35084 39006 35086 39058
rect 35138 39006 35140 39058
rect 35084 38052 35140 39006
rect 35420 39394 35476 39406
rect 35420 39342 35422 39394
rect 35474 39342 35476 39394
rect 35420 39060 35476 39342
rect 37772 39060 37828 39070
rect 35420 39058 35700 39060
rect 35420 39006 35422 39058
rect 35474 39006 35700 39058
rect 35420 39004 35700 39006
rect 35420 38994 35476 39004
rect 35532 38724 35588 38734
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35532 38274 35588 38668
rect 35532 38222 35534 38274
rect 35586 38222 35588 38274
rect 35532 38210 35588 38222
rect 35084 37986 35140 37996
rect 34300 37940 34356 37950
rect 32508 36482 32788 36484
rect 32508 36430 32510 36482
rect 32562 36430 32788 36482
rect 32508 36428 32788 36430
rect 33628 37044 33684 37054
rect 33628 36482 33684 36988
rect 34300 36594 34356 37884
rect 35420 37940 35476 37950
rect 35420 37846 35476 37884
rect 34748 37266 34804 37278
rect 34748 37214 34750 37266
rect 34802 37214 34804 37266
rect 34748 37044 34804 37214
rect 34300 36542 34302 36594
rect 34354 36542 34356 36594
rect 34300 36530 34356 36542
rect 34636 36988 34748 37044
rect 33628 36430 33630 36482
rect 33682 36430 33684 36482
rect 32508 36418 32564 36428
rect 29932 34804 29988 34814
rect 29932 34710 29988 34748
rect 31388 34804 31444 34814
rect 31388 34354 31444 34748
rect 31388 34302 31390 34354
rect 31442 34302 31444 34354
rect 31388 34290 31444 34302
rect 31500 34130 31556 36204
rect 32172 36260 32228 36270
rect 32172 36166 32228 36204
rect 31500 34078 31502 34130
rect 31554 34078 31556 34130
rect 31500 34066 31556 34078
rect 32060 35026 32116 35038
rect 32060 34974 32062 35026
rect 32114 34974 32116 35026
rect 32060 34804 32116 34974
rect 32396 34804 32452 34814
rect 32060 34802 32452 34804
rect 32060 34750 32398 34802
rect 32450 34750 32452 34802
rect 32060 34748 32452 34750
rect 31388 33906 31444 33918
rect 31388 33854 31390 33906
rect 31442 33854 31444 33906
rect 31276 33460 31332 33470
rect 31276 33348 31332 33404
rect 31388 33458 31444 33854
rect 31724 33908 31780 33918
rect 31724 33814 31780 33852
rect 31388 33406 31390 33458
rect 31442 33406 31444 33458
rect 31388 33394 31444 33406
rect 31052 33346 31332 33348
rect 31052 33294 31278 33346
rect 31330 33294 31332 33346
rect 31052 33292 31332 33294
rect 30940 33236 30996 33246
rect 30940 32562 30996 33180
rect 30940 32510 30942 32562
rect 30994 32510 30996 32562
rect 30716 32338 30772 32350
rect 30716 32286 30718 32338
rect 30770 32286 30772 32338
rect 30716 32002 30772 32286
rect 30716 31950 30718 32002
rect 30770 31950 30772 32002
rect 30716 31938 30772 31950
rect 29204 31836 29428 31892
rect 29148 31826 29204 31836
rect 28812 31556 28868 31566
rect 28812 31106 28868 31500
rect 28812 31054 28814 31106
rect 28866 31054 28868 31106
rect 28812 31042 28868 31054
rect 28140 30942 28142 30994
rect 28194 30942 28196 30994
rect 28140 30930 28196 30942
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 29372 28644 29428 31836
rect 30492 31554 30548 31566
rect 30492 31502 30494 31554
rect 30546 31502 30548 31554
rect 30492 30324 30548 31502
rect 30604 31556 30660 31566
rect 30604 31462 30660 31500
rect 30940 30882 30996 32510
rect 31052 32450 31108 33292
rect 31276 33282 31332 33292
rect 31612 33236 31668 33246
rect 31612 33142 31668 33180
rect 31836 33236 31892 33246
rect 32060 33236 32116 34748
rect 32396 34738 32452 34748
rect 32508 34690 32564 34702
rect 32508 34638 32510 34690
rect 32562 34638 32564 34690
rect 32396 34244 32452 34254
rect 32172 34242 32452 34244
rect 32172 34190 32398 34242
rect 32450 34190 32452 34242
rect 32172 34188 32452 34190
rect 32172 33348 32228 34188
rect 32396 34178 32452 34188
rect 32508 34242 32564 34638
rect 32508 34190 32510 34242
rect 32562 34190 32564 34242
rect 32508 34178 32564 34190
rect 32172 33254 32228 33292
rect 32396 33906 32452 33918
rect 32396 33854 32398 33906
rect 32450 33854 32452 33906
rect 32396 33348 32452 33854
rect 32620 33572 32676 36428
rect 33628 36418 33684 36430
rect 33404 34130 33460 34142
rect 33404 34078 33406 34130
rect 33458 34078 33460 34130
rect 33180 33572 33236 33582
rect 32620 33570 33236 33572
rect 32620 33518 33182 33570
rect 33234 33518 33236 33570
rect 32620 33516 33236 33518
rect 33180 33506 33236 33516
rect 33404 33460 33460 34078
rect 33628 33906 33684 33918
rect 33628 33854 33630 33906
rect 33682 33854 33684 33906
rect 33628 33684 33684 33854
rect 33852 33908 33908 33918
rect 33852 33814 33908 33852
rect 33964 33906 34020 33918
rect 33964 33854 33966 33906
rect 34018 33854 34020 33906
rect 33292 33404 33404 33460
rect 32396 33282 32452 33292
rect 32732 33346 32788 33358
rect 32732 33294 32734 33346
rect 32786 33294 32788 33346
rect 31836 33234 32116 33236
rect 31836 33182 31838 33234
rect 31890 33182 32116 33234
rect 31836 33180 32116 33182
rect 31836 33170 31892 33180
rect 32060 33124 32116 33180
rect 32284 33234 32340 33246
rect 32284 33182 32286 33234
rect 32338 33182 32340 33234
rect 32284 33124 32340 33182
rect 32060 33068 32340 33124
rect 32508 33234 32564 33246
rect 32508 33182 32510 33234
rect 32562 33182 32564 33234
rect 31052 32398 31054 32450
rect 31106 32398 31108 32450
rect 31052 32386 31108 32398
rect 31948 33012 32004 33022
rect 31948 32562 32004 32956
rect 31948 32510 31950 32562
rect 32002 32510 32004 32562
rect 31500 31892 31556 31902
rect 31500 31798 31556 31836
rect 30940 30830 30942 30882
rect 30994 30830 30996 30882
rect 30940 30818 30996 30830
rect 31948 30772 32004 32510
rect 32172 32900 32228 32910
rect 32172 32562 32228 32844
rect 32508 32564 32564 33182
rect 32172 32510 32174 32562
rect 32226 32510 32228 32562
rect 32172 31892 32228 32510
rect 32060 31836 32172 31892
rect 32060 30994 32116 31836
rect 32172 31826 32228 31836
rect 32284 32508 32564 32564
rect 32284 31220 32340 32508
rect 32284 31154 32340 31164
rect 32396 32340 32452 32350
rect 32396 31218 32452 32284
rect 32508 32340 32564 32350
rect 32732 32340 32788 33294
rect 32508 32338 32788 32340
rect 32508 32286 32510 32338
rect 32562 32286 32788 32338
rect 32508 32284 32788 32286
rect 32508 32274 32564 32284
rect 32396 31166 32398 31218
rect 32450 31166 32452 31218
rect 32396 31154 32452 31166
rect 32060 30942 32062 30994
rect 32114 30942 32116 30994
rect 32060 30930 32116 30942
rect 32172 30994 32228 31006
rect 32172 30942 32174 30994
rect 32226 30942 32228 30994
rect 32172 30772 32228 30942
rect 32508 30994 32564 31006
rect 32508 30942 32510 30994
rect 32562 30942 32564 30994
rect 32508 30884 32564 30942
rect 32620 30996 32676 32284
rect 33068 31220 33124 31230
rect 33292 31220 33348 33404
rect 33404 33394 33460 33404
rect 33516 33628 33684 33684
rect 33516 32340 33572 33628
rect 33964 33572 34020 33854
rect 33516 32274 33572 32284
rect 33628 33516 34020 33572
rect 33628 31890 33684 33516
rect 33964 33346 34020 33358
rect 33964 33294 33966 33346
rect 34018 33294 34020 33346
rect 33964 32900 34020 33294
rect 34076 33234 34132 33246
rect 34076 33182 34078 33234
rect 34130 33182 34132 33234
rect 34076 33012 34132 33182
rect 34076 32946 34132 32956
rect 33964 32834 34020 32844
rect 34636 32676 34692 36988
rect 34748 36978 34804 36988
rect 35532 37154 35588 37166
rect 35532 37102 35534 37154
rect 35586 37102 35588 37154
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35532 36708 35588 37102
rect 35532 36642 35588 36652
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35420 34356 35476 34366
rect 35644 34356 35700 39004
rect 37100 39058 38164 39060
rect 37100 39006 37774 39058
rect 37826 39006 38164 39058
rect 37100 39004 38164 39006
rect 37100 38946 37156 39004
rect 37772 38994 37828 39004
rect 37100 38894 37102 38946
rect 37154 38894 37156 38946
rect 36988 38724 37044 38762
rect 36988 38658 37044 38668
rect 35756 38052 35812 38062
rect 35756 37958 35812 37996
rect 35980 38052 36036 38062
rect 35980 37958 36036 37996
rect 36988 38050 37044 38062
rect 36988 37998 36990 38050
rect 37042 37998 37044 38050
rect 36428 37828 36484 37838
rect 36988 37828 37044 37998
rect 36428 37826 37044 37828
rect 36428 37774 36430 37826
rect 36482 37774 37044 37826
rect 36428 37772 37044 37774
rect 36428 37762 36484 37772
rect 36428 36932 36484 36942
rect 36428 36594 36484 36876
rect 36428 36542 36430 36594
rect 36482 36542 36484 36594
rect 36428 36530 36484 36542
rect 35420 34354 35644 34356
rect 35420 34302 35422 34354
rect 35474 34302 35644 34354
rect 35420 34300 35644 34302
rect 35420 34290 35476 34300
rect 35644 34262 35700 34300
rect 36204 34356 36260 34366
rect 35084 34242 35140 34254
rect 35084 34190 35086 34242
rect 35138 34190 35140 34242
rect 35084 33908 35140 34190
rect 34748 33460 34804 33470
rect 34748 33366 34804 33404
rect 34972 33348 35028 33358
rect 34972 33254 35028 33292
rect 33628 31838 33630 31890
rect 33682 31838 33684 31890
rect 33628 31826 33684 31838
rect 34412 32674 34692 32676
rect 34412 32622 34638 32674
rect 34690 32622 34692 32674
rect 34412 32620 34692 32622
rect 34412 31778 34468 32620
rect 34636 32610 34692 32620
rect 34412 31726 34414 31778
rect 34466 31726 34468 31778
rect 34412 31714 34468 31726
rect 33068 31218 33348 31220
rect 33068 31166 33070 31218
rect 33122 31166 33348 31218
rect 33068 31164 33348 31166
rect 34300 31220 34356 31230
rect 33068 31154 33124 31164
rect 34300 31126 34356 31164
rect 33964 31106 34020 31118
rect 33964 31054 33966 31106
rect 34018 31054 34020 31106
rect 33404 30996 33460 31006
rect 32620 30994 33460 30996
rect 32620 30942 33406 30994
rect 33458 30942 33460 30994
rect 32620 30940 33460 30942
rect 33404 30930 33460 30940
rect 32508 30818 32564 30828
rect 33628 30884 33684 30894
rect 33964 30884 34020 31054
rect 33684 30828 34020 30884
rect 33628 30790 33684 30828
rect 31948 30716 32340 30772
rect 30492 30258 30548 30268
rect 31388 30324 31444 30334
rect 31388 29650 31444 30268
rect 31388 29598 31390 29650
rect 31442 29598 31444 29650
rect 31388 29586 31444 29598
rect 30156 29204 30212 29214
rect 30156 28754 30212 29148
rect 31276 29204 31332 29214
rect 31612 29204 31668 29214
rect 31276 29110 31332 29148
rect 31500 29202 31668 29204
rect 31500 29150 31614 29202
rect 31666 29150 31668 29202
rect 31500 29148 31668 29150
rect 30156 28702 30158 28754
rect 30210 28702 30212 28754
rect 30156 28690 30212 28702
rect 29372 28550 29428 28588
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 31500 27746 31556 29148
rect 31612 29138 31668 29148
rect 32172 29204 32228 29214
rect 31500 27694 31502 27746
rect 31554 27694 31556 27746
rect 31500 27682 31556 27694
rect 32172 27746 32228 29148
rect 32284 28754 32340 30716
rect 33516 29428 33572 29438
rect 33516 29334 33572 29372
rect 32284 28702 32286 28754
rect 32338 28702 32340 28754
rect 32284 27858 32340 28702
rect 33404 29202 33460 29214
rect 33404 29150 33406 29202
rect 33458 29150 33460 29202
rect 33404 28754 33460 29150
rect 33740 29204 33796 30828
rect 35084 29428 35140 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 36204 33346 36260 34300
rect 36204 33294 36206 33346
rect 36258 33294 36260 33346
rect 36204 33282 36260 33294
rect 35644 33236 35700 33246
rect 35644 33234 35812 33236
rect 35644 33182 35646 33234
rect 35698 33182 35812 33234
rect 35644 33180 35812 33182
rect 35644 33170 35700 33180
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35644 30994 35700 31006
rect 35644 30942 35646 30994
rect 35698 30942 35700 30994
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35644 30436 35700 30942
rect 35756 30770 35812 33180
rect 35980 33124 36036 33134
rect 35980 33030 36036 33068
rect 35980 31668 36036 31678
rect 35868 31612 35980 31668
rect 35868 31218 35924 31612
rect 35980 31602 36036 31612
rect 35868 31166 35870 31218
rect 35922 31166 35924 31218
rect 35868 31154 35924 31166
rect 36092 31556 36148 31566
rect 36092 31218 36148 31500
rect 36092 31166 36094 31218
rect 36146 31166 36148 31218
rect 36092 31154 36148 31166
rect 36316 31108 36372 31118
rect 36316 31014 36372 31052
rect 36540 30772 36596 37772
rect 36988 36708 37044 36718
rect 36988 36614 37044 36652
rect 37100 36370 37156 38894
rect 37996 38834 38052 38846
rect 37996 38782 37998 38834
rect 38050 38782 38052 38834
rect 37996 38668 38052 38782
rect 37324 38610 37380 38622
rect 37324 38558 37326 38610
rect 37378 38558 37380 38610
rect 37324 36932 37380 38558
rect 37324 36866 37380 36876
rect 37660 38612 38052 38668
rect 37660 37154 37716 38612
rect 37996 37268 38052 37278
rect 38108 37268 38164 39004
rect 39340 38668 39396 39678
rect 39452 38834 39508 38846
rect 39452 38782 39454 38834
rect 39506 38782 39508 38834
rect 39452 38668 39508 38782
rect 39340 38612 39508 38668
rect 39228 38164 39284 38174
rect 38556 38052 38612 38062
rect 38556 37490 38612 37996
rect 38556 37438 38558 37490
rect 38610 37438 38612 37490
rect 38556 37426 38612 37438
rect 37996 37266 38164 37268
rect 37996 37214 37998 37266
rect 38050 37214 38164 37266
rect 37996 37212 38164 37214
rect 37996 37202 38052 37212
rect 37660 37102 37662 37154
rect 37714 37102 37716 37154
rect 37660 36596 37716 37102
rect 37996 37044 38052 37054
rect 37996 36706 38052 36988
rect 37996 36654 37998 36706
rect 38050 36654 38052 36706
rect 37996 36642 38052 36654
rect 38108 36706 38164 37212
rect 38220 37042 38276 37054
rect 38220 36990 38222 37042
rect 38274 36990 38276 37042
rect 38220 36932 38276 36990
rect 38276 36876 38388 36932
rect 38220 36866 38276 36876
rect 38108 36654 38110 36706
rect 38162 36654 38164 36706
rect 38108 36642 38164 36654
rect 38332 36706 38388 36876
rect 38332 36654 38334 36706
rect 38386 36654 38388 36706
rect 38332 36642 38388 36654
rect 39116 36820 39172 36830
rect 37660 36530 37716 36540
rect 38892 36596 38948 36606
rect 38892 36502 38948 36540
rect 38444 36484 38500 36494
rect 37996 36482 38500 36484
rect 37996 36430 38446 36482
rect 38498 36430 38500 36482
rect 37996 36428 38500 36430
rect 37100 36318 37102 36370
rect 37154 36318 37156 36370
rect 37100 36306 37156 36318
rect 37324 36372 37380 36382
rect 37324 36278 37380 36316
rect 37100 34356 37156 34366
rect 37100 34262 37156 34300
rect 37436 34244 37492 34254
rect 37436 34150 37492 34188
rect 37436 33458 37492 33470
rect 37436 33406 37438 33458
rect 37490 33406 37492 33458
rect 36988 31778 37044 31790
rect 36988 31726 36990 31778
rect 37042 31726 37044 31778
rect 36764 30996 36820 31006
rect 36764 30902 36820 30940
rect 35756 30718 35758 30770
rect 35810 30718 35812 30770
rect 35756 30706 35812 30718
rect 36316 30716 36596 30772
rect 36204 30436 36260 30446
rect 35532 30380 36148 30436
rect 35196 29428 35252 29438
rect 35084 29372 35196 29428
rect 35196 29334 35252 29372
rect 33740 29110 33796 29148
rect 33852 29202 33908 29214
rect 35084 29204 35140 29214
rect 33852 29150 33854 29202
rect 33906 29150 33908 29202
rect 33852 28868 33908 29150
rect 33852 28802 33908 28812
rect 34748 29202 35140 29204
rect 34748 29150 35086 29202
rect 35138 29150 35140 29202
rect 34748 29148 35140 29150
rect 33404 28702 33406 28754
rect 33458 28702 33460 28754
rect 33404 28690 33460 28702
rect 32620 28644 32676 28654
rect 32620 28550 32676 28588
rect 33964 28644 34020 28654
rect 32284 27806 32286 27858
rect 32338 27806 32340 27858
rect 32284 27794 32340 27806
rect 33964 27858 34020 28588
rect 34748 27970 34804 29148
rect 35084 29138 35140 29148
rect 35420 29204 35476 29242
rect 35420 29138 35476 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35532 28756 35588 30380
rect 36092 30322 36148 30380
rect 36092 30270 36094 30322
rect 36146 30270 36148 30322
rect 36092 30258 36148 30270
rect 36204 30210 36260 30380
rect 36204 30158 36206 30210
rect 36258 30158 36260 30210
rect 36204 30146 36260 30158
rect 36204 29652 36260 29662
rect 35644 29426 35700 29438
rect 35644 29374 35646 29426
rect 35698 29374 35700 29426
rect 35644 29204 35700 29374
rect 36204 29426 36260 29596
rect 36204 29374 36206 29426
rect 36258 29374 36260 29426
rect 36204 29362 36260 29374
rect 36092 29204 36148 29214
rect 35644 29202 36148 29204
rect 35644 29150 36094 29202
rect 36146 29150 36148 29202
rect 35644 29148 36148 29150
rect 35980 28868 36036 28878
rect 36092 28868 36148 29148
rect 36204 28868 36260 28878
rect 36092 28866 36260 28868
rect 36092 28814 36206 28866
rect 36258 28814 36260 28866
rect 36092 28812 36260 28814
rect 35532 28754 35924 28756
rect 35532 28702 35534 28754
rect 35586 28702 35924 28754
rect 35532 28700 35924 28702
rect 35532 28690 35588 28700
rect 35868 28642 35924 28700
rect 35980 28754 36036 28812
rect 36204 28802 36260 28812
rect 35980 28702 35982 28754
rect 36034 28702 36036 28754
rect 35980 28690 36036 28702
rect 35868 28590 35870 28642
rect 35922 28590 35924 28642
rect 35868 28578 35924 28590
rect 34748 27918 34750 27970
rect 34802 27918 34804 27970
rect 34748 27906 34804 27918
rect 33964 27806 33966 27858
rect 34018 27806 34020 27858
rect 33964 27794 34020 27806
rect 32172 27694 32174 27746
rect 32226 27694 32228 27746
rect 32172 27682 32228 27694
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 36316 20188 36372 30716
rect 36988 30436 37044 31726
rect 36988 30370 37044 30380
rect 37100 31668 37156 31678
rect 37100 29652 37156 31612
rect 37212 31554 37268 31566
rect 37212 31502 37214 31554
rect 37266 31502 37268 31554
rect 37212 31220 37268 31502
rect 37212 31154 37268 31164
rect 37436 31106 37492 33406
rect 37772 33234 37828 33246
rect 37772 33182 37774 33234
rect 37826 33182 37828 33234
rect 37436 31054 37438 31106
rect 37490 31054 37492 31106
rect 37436 31042 37492 31054
rect 37548 33124 37604 33134
rect 37548 30324 37604 33068
rect 37548 29652 37604 30268
rect 37772 30210 37828 33182
rect 37772 30158 37774 30210
rect 37826 30158 37828 30210
rect 37772 30146 37828 30158
rect 37996 31778 38052 36428
rect 38444 36418 38500 36428
rect 39116 36482 39172 36764
rect 39116 36430 39118 36482
rect 39170 36430 39172 36482
rect 39116 36418 39172 36430
rect 38668 34916 38724 34926
rect 38668 34822 38724 34860
rect 38892 34244 38948 34254
rect 38332 33348 38388 33358
rect 38332 32562 38388 33292
rect 38332 32510 38334 32562
rect 38386 32510 38388 32562
rect 38332 32498 38388 32510
rect 38556 32004 38612 32014
rect 38556 31780 38612 31948
rect 37996 31726 37998 31778
rect 38050 31726 38052 31778
rect 37772 29652 37828 29662
rect 37548 29596 37772 29652
rect 37100 29558 37156 29596
rect 37772 29586 37828 29596
rect 37884 29652 37940 29662
rect 37996 29652 38052 31726
rect 37884 29650 38052 29652
rect 37884 29598 37886 29650
rect 37938 29598 38052 29650
rect 37884 29596 38052 29598
rect 38108 31724 38612 31780
rect 36652 29428 36708 29438
rect 36652 29334 36708 29372
rect 36428 29316 36484 29326
rect 36428 29222 36484 29260
rect 36988 29314 37044 29326
rect 36988 29262 36990 29314
rect 37042 29262 37044 29314
rect 36540 29204 36596 29214
rect 36540 27300 36596 29148
rect 36876 27748 36932 27758
rect 36988 27748 37044 29262
rect 37884 29316 37940 29596
rect 38108 29540 38164 31724
rect 38556 31666 38612 31724
rect 38556 31614 38558 31666
rect 38610 31614 38612 31666
rect 38556 31602 38612 31614
rect 38444 31556 38500 31566
rect 38444 30210 38500 31500
rect 38892 30436 38948 34188
rect 39228 33348 39284 38108
rect 39340 36372 39396 38612
rect 39564 38164 39620 41132
rect 39564 38070 39620 38108
rect 39676 37492 39732 41694
rect 39900 41300 39956 43262
rect 40348 43092 40404 43598
rect 40348 43026 40404 43036
rect 42028 43540 42084 44268
rect 43372 44996 43428 45006
rect 42140 44212 42196 44222
rect 42140 44118 42196 44156
rect 43372 43650 43428 44940
rect 44268 44436 44324 44446
rect 44828 44436 44884 44446
rect 44268 44434 44884 44436
rect 44268 44382 44270 44434
rect 44322 44382 44830 44434
rect 44882 44382 44884 44434
rect 44268 44380 44884 44382
rect 45052 44436 45108 48972
rect 45612 48914 45668 48926
rect 45612 48862 45614 48914
rect 45666 48862 45668 48914
rect 45612 48466 45668 48862
rect 45612 48414 45614 48466
rect 45666 48414 45668 48466
rect 45612 48402 45668 48414
rect 47628 48468 47684 48478
rect 47628 48374 47684 48412
rect 45836 48354 45892 48366
rect 45836 48302 45838 48354
rect 45890 48302 45892 48354
rect 45500 47348 45556 47358
rect 45164 47346 45556 47348
rect 45164 47294 45502 47346
rect 45554 47294 45556 47346
rect 45164 47292 45556 47294
rect 45164 46562 45220 47292
rect 45500 47282 45556 47292
rect 45612 47234 45668 47246
rect 45612 47182 45614 47234
rect 45666 47182 45668 47234
rect 45612 47124 45668 47182
rect 45164 46510 45166 46562
rect 45218 46510 45220 46562
rect 45164 46498 45220 46510
rect 45500 47068 45668 47124
rect 45836 47124 45892 48302
rect 47740 48356 47796 48366
rect 47740 48262 47796 48300
rect 45948 48244 46004 48254
rect 47404 48244 47460 48254
rect 45948 48242 46452 48244
rect 45948 48190 45950 48242
rect 46002 48190 46452 48242
rect 45948 48188 46452 48190
rect 45948 48178 46004 48188
rect 46284 48020 46340 48030
rect 46284 47346 46340 47964
rect 46396 47458 46452 48188
rect 47292 48242 47460 48244
rect 47292 48190 47406 48242
rect 47458 48190 47460 48242
rect 47292 48188 47460 48190
rect 46732 47516 47124 47572
rect 46732 47460 46788 47516
rect 46396 47406 46398 47458
rect 46450 47406 46452 47458
rect 46396 47394 46452 47406
rect 46508 47458 46788 47460
rect 46508 47406 46734 47458
rect 46786 47406 46788 47458
rect 46508 47404 46788 47406
rect 46284 47294 46286 47346
rect 46338 47294 46340 47346
rect 46284 47236 46340 47294
rect 46284 47170 46340 47180
rect 45500 46676 45556 47068
rect 45836 47058 45892 47068
rect 46508 47012 46564 47404
rect 46732 47394 46788 47404
rect 46844 47348 46900 47358
rect 46620 47236 46676 47246
rect 46620 47142 46676 47180
rect 46284 46956 46564 47012
rect 46732 47124 46788 47134
rect 46172 46676 46228 46686
rect 46284 46676 46340 46956
rect 46620 46900 46676 46910
rect 46732 46900 46788 47068
rect 46620 46898 46788 46900
rect 46620 46846 46622 46898
rect 46674 46846 46788 46898
rect 46620 46844 46788 46846
rect 46620 46834 46676 46844
rect 46844 46786 46900 47292
rect 47068 47346 47124 47516
rect 47068 47294 47070 47346
rect 47122 47294 47124 47346
rect 47068 47282 47124 47294
rect 46844 46734 46846 46786
rect 46898 46734 46900 46786
rect 46844 46722 46900 46734
rect 45276 45220 45332 45230
rect 45052 44380 45220 44436
rect 44268 44370 44324 44380
rect 44828 44370 44884 44380
rect 44940 44100 44996 44110
rect 44940 44006 44996 44044
rect 43372 43598 43374 43650
rect 43426 43598 43428 43650
rect 43372 43586 43428 43598
rect 42588 43540 42644 43550
rect 42028 43538 42644 43540
rect 42028 43486 42590 43538
rect 42642 43486 42644 43538
rect 42028 43484 42644 43486
rect 42028 42866 42084 43484
rect 42588 43474 42644 43484
rect 42028 42814 42030 42866
rect 42082 42814 42084 42866
rect 40796 41972 40852 41982
rect 40796 41878 40852 41916
rect 41132 41972 41188 41982
rect 41132 41878 41188 41916
rect 41356 41970 41412 41982
rect 41356 41918 41358 41970
rect 41410 41918 41412 41970
rect 39900 41234 39956 41244
rect 41020 41858 41076 41870
rect 41020 41806 41022 41858
rect 41074 41806 41076 41858
rect 41020 40516 41076 41806
rect 41244 41300 41300 41310
rect 41244 41206 41300 41244
rect 41020 40450 41076 40460
rect 41132 40068 41188 40078
rect 41356 40068 41412 41918
rect 41468 41188 41524 41198
rect 41468 40626 41524 41132
rect 42028 41186 42084 42814
rect 44604 42196 44660 42206
rect 45164 42196 45220 44380
rect 45276 44322 45332 45164
rect 45276 44270 45278 44322
rect 45330 44270 45332 44322
rect 45276 44258 45332 44270
rect 45388 44212 45444 44222
rect 45388 44118 45444 44156
rect 45500 43988 45556 46620
rect 46060 46674 46340 46676
rect 46060 46622 46174 46674
rect 46226 46622 46340 46674
rect 46060 46620 46340 46622
rect 46396 46676 46452 46686
rect 46060 45220 46116 46620
rect 46172 46610 46228 46620
rect 46396 46582 46452 46620
rect 46508 46564 46564 46574
rect 46508 46470 46564 46508
rect 47180 46116 47236 46126
rect 47292 46116 47348 48188
rect 47404 48178 47460 48188
rect 47516 48130 47572 48142
rect 47516 48078 47518 48130
rect 47570 48078 47572 48130
rect 47404 47234 47460 47246
rect 47404 47182 47406 47234
rect 47458 47182 47460 47234
rect 47404 46900 47460 47182
rect 47516 47124 47572 48078
rect 47852 48020 47908 49084
rect 49532 49140 49588 55412
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 78204 50370 78260 50382
rect 78204 50318 78206 50370
rect 78258 50318 78260 50370
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 78204 49812 78260 50318
rect 78204 49746 78260 49756
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 49532 49074 49588 49084
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 48748 48468 48804 48478
rect 48188 48244 48244 48254
rect 48188 48242 48580 48244
rect 48188 48190 48190 48242
rect 48242 48190 48580 48242
rect 48188 48188 48580 48190
rect 48188 48178 48244 48188
rect 47852 47954 47908 47964
rect 47852 47458 47908 47470
rect 47852 47406 47854 47458
rect 47906 47406 47908 47458
rect 47740 47348 47796 47358
rect 47740 47254 47796 47292
rect 47852 47124 47908 47406
rect 47516 47058 47572 47068
rect 47628 47068 47908 47124
rect 48076 47458 48132 47470
rect 48076 47406 48078 47458
rect 48130 47406 48132 47458
rect 47628 47012 47684 47068
rect 47628 46900 47684 46956
rect 47404 46844 47684 46900
rect 47404 46676 47460 46686
rect 47460 46620 47572 46676
rect 47404 46610 47460 46620
rect 47516 46452 47572 46620
rect 47628 46674 47684 46686
rect 47628 46622 47630 46674
rect 47682 46622 47684 46674
rect 47628 46564 47684 46622
rect 47740 46676 47796 46686
rect 47740 46582 47796 46620
rect 47964 46674 48020 46686
rect 47964 46622 47966 46674
rect 48018 46622 48020 46674
rect 47628 46498 47684 46508
rect 47964 46452 48020 46622
rect 47516 46340 47572 46396
rect 47740 46396 48020 46452
rect 48076 46452 48132 47406
rect 48188 47460 48244 47470
rect 48188 46786 48244 47404
rect 48300 47458 48356 47470
rect 48300 47406 48302 47458
rect 48354 47406 48356 47458
rect 48300 47236 48356 47406
rect 48300 47170 48356 47180
rect 48188 46734 48190 46786
rect 48242 46734 48244 46786
rect 48188 46722 48244 46734
rect 48300 46788 48356 46798
rect 48300 46694 48356 46732
rect 48524 46676 48580 48188
rect 48748 47572 48804 48412
rect 49756 48356 49812 48366
rect 49084 48244 49140 48254
rect 49084 48150 49140 48188
rect 49532 48132 49588 48142
rect 49532 48038 49588 48076
rect 49420 48020 49476 48030
rect 48748 47506 48804 47516
rect 49196 48018 49476 48020
rect 49196 47966 49422 48018
rect 49474 47966 49476 48018
rect 49196 47964 49476 47966
rect 48860 47458 48916 47470
rect 48860 47406 48862 47458
rect 48914 47406 48916 47458
rect 48636 47236 48692 47246
rect 48636 47142 48692 47180
rect 48860 46900 48916 47406
rect 48076 46396 48468 46452
rect 47516 46284 47684 46340
rect 47516 46116 47572 46126
rect 47292 46114 47572 46116
rect 47292 46062 47518 46114
rect 47570 46062 47572 46114
rect 47292 46060 47572 46062
rect 47180 46022 47236 46060
rect 47516 46050 47572 46060
rect 46844 46004 46900 46014
rect 46060 45126 46116 45164
rect 46172 46002 46900 46004
rect 46172 45950 46846 46002
rect 46898 45950 46900 46002
rect 46172 45948 46900 45950
rect 45836 45108 45892 45118
rect 45836 45014 45892 45052
rect 45948 44996 46004 45006
rect 45948 44902 46004 44940
rect 46172 44772 46228 45948
rect 46844 45938 46900 45948
rect 47628 46002 47684 46284
rect 47628 45950 47630 46002
rect 47682 45950 47684 46002
rect 47628 45938 47684 45950
rect 47740 45780 47796 46396
rect 48412 46114 48468 46396
rect 48412 46062 48414 46114
rect 48466 46062 48468 46114
rect 48412 46050 48468 46062
rect 48300 45892 48356 45902
rect 48524 45892 48580 46620
rect 48300 45890 48580 45892
rect 48300 45838 48302 45890
rect 48354 45838 48580 45890
rect 48300 45836 48580 45838
rect 48636 46844 48916 46900
rect 48972 47458 49028 47470
rect 48972 47406 48974 47458
rect 49026 47406 49028 47458
rect 48636 46564 48692 46844
rect 48748 46676 48804 46686
rect 48748 46582 48804 46620
rect 48636 45890 48692 46508
rect 48860 46452 48916 46462
rect 48860 46358 48916 46396
rect 48972 45892 49028 47406
rect 49196 47460 49252 47964
rect 49420 47954 49476 47964
rect 49196 47366 49252 47404
rect 49420 47572 49476 47582
rect 49756 47572 49812 48300
rect 49980 48244 50036 48254
rect 49980 48132 50036 48188
rect 50876 48244 50932 48254
rect 50876 48242 51380 48244
rect 50876 48190 50878 48242
rect 50930 48190 51380 48242
rect 50876 48188 51380 48190
rect 50876 48178 50932 48188
rect 50540 48132 50596 48142
rect 49980 48130 50372 48132
rect 49980 48078 49982 48130
rect 50034 48078 50372 48130
rect 49980 48076 50372 48078
rect 49980 48066 50036 48076
rect 49756 47516 50260 47572
rect 49420 47460 49476 47516
rect 49420 47458 49700 47460
rect 49420 47406 49422 47458
rect 49474 47406 49700 47458
rect 49420 47404 49700 47406
rect 49420 47394 49476 47404
rect 49420 46900 49476 46910
rect 49084 46788 49140 46798
rect 49420 46788 49476 46844
rect 49084 46694 49140 46732
rect 49196 46786 49476 46788
rect 49196 46734 49422 46786
rect 49474 46734 49476 46786
rect 49196 46732 49476 46734
rect 48636 45838 48638 45890
rect 48690 45838 48692 45890
rect 48300 45826 48356 45836
rect 47964 45780 48020 45790
rect 47740 45778 48020 45780
rect 47740 45726 47966 45778
rect 48018 45726 48020 45778
rect 47740 45724 48020 45726
rect 46956 45666 47012 45678
rect 46956 45614 46958 45666
rect 47010 45614 47012 45666
rect 46956 45556 47012 45614
rect 45836 44716 46228 44772
rect 46396 45106 46452 45118
rect 46396 45054 46398 45106
rect 46450 45054 46452 45106
rect 45836 44322 45892 44716
rect 46396 44546 46452 45054
rect 46396 44494 46398 44546
rect 46450 44494 46452 44546
rect 46396 44482 46452 44494
rect 45836 44270 45838 44322
rect 45890 44270 45892 44322
rect 45836 44258 45892 44270
rect 46508 44324 46564 44334
rect 46956 44324 47012 45500
rect 47964 45332 48020 45724
rect 48636 45780 48692 45838
rect 48636 45714 48692 45724
rect 48748 45836 49028 45892
rect 49084 45892 49140 45902
rect 49196 45892 49252 46732
rect 49420 46722 49476 46732
rect 49644 46786 49700 47404
rect 49644 46734 49646 46786
rect 49698 46734 49700 46786
rect 49644 46564 49700 46734
rect 49868 47346 49924 47358
rect 49868 47294 49870 47346
rect 49922 47294 49924 47346
rect 49084 45890 49252 45892
rect 49084 45838 49086 45890
rect 49138 45838 49252 45890
rect 49084 45836 49252 45838
rect 49308 46508 49700 46564
rect 49756 46562 49812 46574
rect 49756 46510 49758 46562
rect 49810 46510 49812 46562
rect 48076 45668 48132 45678
rect 48076 45574 48132 45612
rect 48748 45444 48804 45836
rect 49084 45826 49140 45836
rect 49308 45778 49364 46508
rect 49308 45726 49310 45778
rect 49362 45726 49364 45778
rect 49308 45714 49364 45726
rect 49420 46228 49476 46238
rect 49420 46002 49476 46172
rect 49756 46116 49812 46510
rect 49868 46452 49924 47294
rect 49980 47234 50036 47246
rect 49980 47182 49982 47234
rect 50034 47182 50036 47234
rect 49980 46676 50036 47182
rect 50092 46786 50148 47516
rect 50204 47458 50260 47516
rect 50204 47406 50206 47458
rect 50258 47406 50260 47458
rect 50204 47394 50260 47406
rect 50316 47236 50372 48076
rect 50540 47684 50596 48076
rect 51100 47684 51156 47694
rect 50540 47618 50596 47628
rect 50988 47628 51100 47684
rect 50540 47236 50596 47246
rect 50316 47234 50596 47236
rect 50316 47182 50542 47234
rect 50594 47182 50596 47234
rect 50316 47180 50596 47182
rect 50092 46734 50094 46786
rect 50146 46734 50148 46786
rect 50092 46722 50148 46734
rect 50204 47012 50260 47022
rect 50204 46898 50260 46956
rect 50204 46846 50206 46898
rect 50258 46846 50260 46898
rect 49980 46610 50036 46620
rect 49924 46396 50036 46452
rect 49868 46386 49924 46396
rect 49756 46050 49812 46060
rect 49420 45950 49422 46002
rect 49474 45950 49476 46002
rect 47068 45108 47124 45118
rect 47068 45014 47124 45052
rect 47964 45106 48020 45276
rect 47964 45054 47966 45106
rect 48018 45054 48020 45106
rect 47964 45042 48020 45054
rect 48636 45388 48804 45444
rect 49420 45668 49476 45950
rect 47852 44996 47908 45006
rect 47852 44902 47908 44940
rect 48636 44996 48692 45388
rect 48860 45332 48916 45342
rect 48860 45238 48916 45276
rect 49420 45330 49476 45612
rect 49868 45666 49924 45678
rect 49868 45614 49870 45666
rect 49922 45614 49924 45666
rect 49868 45556 49924 45614
rect 49868 45490 49924 45500
rect 49420 45278 49422 45330
rect 49474 45278 49476 45330
rect 49420 45266 49476 45278
rect 49980 45330 50036 46396
rect 50204 45890 50260 46846
rect 50316 46788 50372 46798
rect 50316 46694 50372 46732
rect 50204 45838 50206 45890
rect 50258 45838 50260 45890
rect 50204 45826 50260 45838
rect 50428 45892 50484 47180
rect 50540 47170 50596 47180
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50876 46676 50932 46686
rect 50876 46004 50932 46620
rect 50988 46228 51044 47628
rect 51100 47618 51156 47628
rect 51100 46900 51156 46910
rect 51100 46806 51156 46844
rect 50988 46004 51044 46172
rect 51100 46004 51156 46014
rect 50988 46002 51156 46004
rect 50988 45950 51102 46002
rect 51154 45950 51156 46002
rect 50988 45948 51156 45950
rect 50876 45938 50932 45948
rect 51100 45938 51156 45948
rect 50652 45892 50708 45902
rect 50428 45836 50652 45892
rect 49980 45278 49982 45330
rect 50034 45278 50036 45330
rect 49980 45266 50036 45278
rect 50316 45780 50372 45790
rect 50204 45218 50260 45230
rect 50204 45166 50206 45218
rect 50258 45166 50260 45218
rect 48636 44930 48692 44940
rect 49868 45106 49924 45118
rect 49868 45054 49870 45106
rect 49922 45054 49924 45106
rect 49868 44548 49924 45054
rect 49868 44454 49924 44492
rect 46508 44322 47012 44324
rect 46508 44270 46510 44322
rect 46562 44270 47012 44322
rect 46508 44268 47012 44270
rect 46508 44258 46564 44268
rect 45612 44212 45668 44222
rect 45612 44210 45780 44212
rect 45612 44158 45614 44210
rect 45666 44158 45780 44210
rect 45612 44156 45780 44158
rect 45612 44146 45668 44156
rect 44604 42194 45220 42196
rect 44604 42142 44606 42194
rect 44658 42142 45220 42194
rect 44604 42140 45220 42142
rect 43036 41300 43092 41310
rect 42028 41134 42030 41186
rect 42082 41134 42084 41186
rect 41468 40574 41470 40626
rect 41522 40574 41524 40626
rect 41468 40562 41524 40574
rect 41692 41076 41748 41086
rect 41692 40626 41748 41020
rect 42028 40852 42084 41134
rect 42252 41188 42308 41198
rect 42084 40796 42196 40852
rect 42028 40786 42084 40796
rect 41692 40574 41694 40626
rect 41746 40574 41748 40626
rect 41692 40562 41748 40574
rect 41188 40012 41412 40068
rect 42028 40178 42084 40190
rect 42028 40126 42030 40178
rect 42082 40126 42084 40178
rect 41132 38946 41188 40012
rect 42028 39620 42084 40126
rect 41468 39508 41524 39518
rect 41132 38894 41134 38946
rect 41186 38894 41188 38946
rect 40348 38836 40404 38846
rect 40908 38836 40964 38846
rect 40348 38834 40964 38836
rect 40348 38782 40350 38834
rect 40402 38782 40910 38834
rect 40962 38782 40964 38834
rect 40348 38780 40964 38782
rect 40348 38770 40404 38780
rect 40908 38770 40964 38780
rect 41132 38836 41188 38894
rect 41132 38770 41188 38780
rect 41244 39506 41524 39508
rect 41244 39454 41470 39506
rect 41522 39454 41524 39506
rect 41244 39452 41524 39454
rect 39788 38722 39844 38734
rect 39788 38670 39790 38722
rect 39842 38670 39844 38722
rect 39788 38052 39844 38670
rect 41244 38722 41300 39452
rect 41468 39442 41524 39452
rect 41244 38670 41246 38722
rect 41298 38670 41300 38722
rect 41244 38658 41300 38670
rect 42028 38724 42084 39564
rect 42140 39618 42196 40796
rect 42252 40514 42308 41132
rect 42812 41188 42868 41198
rect 42812 41094 42868 41132
rect 43036 41074 43092 41244
rect 44156 41300 44212 41310
rect 43484 41188 43540 41198
rect 43484 41094 43540 41132
rect 44156 41186 44212 41244
rect 44156 41134 44158 41186
rect 44210 41134 44212 41186
rect 44156 41122 44212 41134
rect 43820 41076 43876 41086
rect 43036 41022 43038 41074
rect 43090 41022 43092 41074
rect 43036 41010 43092 41022
rect 43596 41074 43876 41076
rect 43596 41022 43822 41074
rect 43874 41022 43876 41074
rect 43596 41020 43876 41022
rect 43372 40964 43428 40974
rect 42252 40462 42254 40514
rect 42306 40462 42308 40514
rect 42252 40450 42308 40462
rect 42700 40852 42756 40862
rect 42700 40402 42756 40796
rect 43372 40514 43428 40908
rect 43372 40462 43374 40514
rect 43426 40462 43428 40514
rect 43372 40450 43428 40462
rect 42700 40350 42702 40402
rect 42754 40350 42756 40402
rect 42700 40338 42756 40350
rect 43596 39842 43652 41020
rect 43820 41010 43876 41020
rect 43932 40964 43988 40974
rect 43932 40870 43988 40908
rect 43596 39790 43598 39842
rect 43650 39790 43652 39842
rect 43596 39778 43652 39790
rect 42140 39566 42142 39618
rect 42194 39566 42196 39618
rect 42140 39554 42196 39566
rect 42924 39730 42980 39742
rect 42924 39678 42926 39730
rect 42978 39678 42980 39730
rect 42924 39620 42980 39678
rect 42924 39554 42980 39564
rect 43260 39620 43316 39630
rect 43260 39526 43316 39564
rect 44604 39620 44660 42140
rect 44940 41972 44996 41982
rect 45164 41972 45220 42140
rect 45388 43932 45556 43988
rect 45724 44100 45780 44156
rect 49756 44210 49812 44222
rect 49756 44158 49758 44210
rect 49810 44158 49812 44210
rect 45276 41972 45332 41982
rect 45164 41970 45332 41972
rect 45164 41918 45278 41970
rect 45330 41918 45332 41970
rect 45164 41916 45332 41918
rect 44940 41878 44996 41916
rect 45276 41860 45332 41916
rect 45276 41794 45332 41804
rect 45388 40068 45444 43932
rect 45500 43426 45556 43438
rect 45500 43374 45502 43426
rect 45554 43374 45556 43426
rect 45500 42980 45556 43374
rect 45500 42914 45556 42924
rect 45612 42530 45668 42542
rect 45612 42478 45614 42530
rect 45666 42478 45668 42530
rect 45612 41972 45668 42478
rect 45612 41906 45668 41916
rect 45612 41412 45668 41422
rect 45724 41412 45780 44044
rect 46396 44098 46452 44110
rect 46396 44046 46398 44098
rect 46450 44046 46452 44098
rect 46284 43426 46340 43438
rect 46284 43374 46286 43426
rect 46338 43374 46340 43426
rect 45948 42756 46004 42766
rect 46284 42756 46340 43374
rect 46396 42980 46452 44046
rect 49756 43764 49812 44158
rect 49756 43698 49812 43708
rect 50204 44100 50260 45166
rect 50316 44546 50372 45724
rect 50428 45332 50484 45836
rect 50652 45798 50708 45836
rect 51324 45556 51380 48188
rect 75628 48242 75684 48254
rect 75628 48190 75630 48242
rect 75682 48190 75684 48242
rect 51548 48130 51604 48142
rect 51548 48078 51550 48130
rect 51602 48078 51604 48130
rect 51548 47570 51604 48078
rect 51548 47518 51550 47570
rect 51602 47518 51604 47570
rect 51548 47506 51604 47518
rect 53676 48130 53732 48142
rect 53676 48078 53678 48130
rect 53730 48078 53732 48130
rect 51884 47458 51940 47470
rect 51884 47406 51886 47458
rect 51938 47406 51940 47458
rect 51436 47346 51492 47358
rect 51436 47294 51438 47346
rect 51490 47294 51492 47346
rect 51436 46900 51492 47294
rect 51772 47348 51828 47358
rect 51772 47254 51828 47292
rect 51436 46834 51492 46844
rect 51884 46788 51940 47406
rect 52780 47458 52836 47470
rect 52780 47406 52782 47458
rect 52834 47406 52836 47458
rect 52668 47348 52724 47358
rect 52780 47348 52836 47406
rect 52892 47348 52948 47358
rect 52780 47292 52892 47348
rect 52668 47254 52724 47292
rect 52892 47282 52948 47292
rect 53340 47348 53396 47358
rect 53340 47254 53396 47292
rect 53676 47348 53732 48078
rect 75404 48132 75460 48142
rect 75628 48132 75684 48190
rect 75404 48130 75684 48132
rect 75404 48078 75406 48130
rect 75458 48078 75684 48130
rect 75404 48076 75684 48078
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 53676 47282 53732 47292
rect 75404 47348 75460 48076
rect 77980 48018 78036 48030
rect 77980 47966 77982 48018
rect 78034 47966 78036 48018
rect 77980 47796 78036 47966
rect 77980 47730 78036 47740
rect 75404 47282 75460 47292
rect 77868 47684 77924 47694
rect 77868 47346 77924 47628
rect 77868 47294 77870 47346
rect 77922 47294 77924 47346
rect 77868 47282 77924 47294
rect 77644 47234 77700 47246
rect 77644 47182 77646 47234
rect 77698 47182 77700 47234
rect 77644 47124 77700 47182
rect 77644 47058 77700 47068
rect 78204 47234 78260 47246
rect 78204 47182 78206 47234
rect 78258 47182 78260 47234
rect 78204 47124 78260 47182
rect 78204 47058 78260 47068
rect 51772 46732 51884 46788
rect 51436 45780 51492 45790
rect 51436 45686 51492 45724
rect 51548 45666 51604 45678
rect 51548 45614 51550 45666
rect 51602 45614 51604 45666
rect 50556 45500 50820 45510
rect 51324 45500 51492 45556
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50428 45266 50484 45276
rect 50652 45220 50708 45230
rect 50652 45126 50708 45164
rect 51436 45108 51492 45500
rect 50764 45106 51492 45108
rect 50764 45054 51438 45106
rect 51490 45054 51492 45106
rect 50764 45052 51492 45054
rect 50316 44494 50318 44546
rect 50370 44494 50372 44546
rect 50316 44482 50372 44494
rect 50428 44548 50484 44558
rect 50428 44322 50484 44492
rect 50428 44270 50430 44322
rect 50482 44270 50484 44322
rect 50428 44258 50484 44270
rect 50316 44100 50372 44110
rect 50764 44100 50820 45052
rect 51436 45042 51492 45052
rect 51548 45108 51604 45614
rect 51660 45666 51716 45678
rect 51660 45614 51662 45666
rect 51714 45614 51716 45666
rect 51660 45556 51716 45614
rect 51660 45490 51716 45500
rect 51548 45042 51604 45052
rect 50204 44098 50372 44100
rect 50204 44046 50318 44098
rect 50370 44046 50372 44098
rect 50204 44044 50372 44046
rect 48188 43652 48244 43662
rect 46396 42914 46452 42924
rect 47404 42980 47460 42990
rect 47404 42886 47460 42924
rect 46844 42756 46900 42766
rect 45948 42754 46900 42756
rect 45948 42702 45950 42754
rect 46002 42702 46846 42754
rect 46898 42702 46900 42754
rect 45948 42700 46900 42702
rect 45948 42690 46004 42700
rect 46284 42532 46340 42542
rect 46172 42530 46340 42532
rect 46172 42478 46286 42530
rect 46338 42478 46340 42530
rect 46172 42476 46340 42478
rect 46060 41860 46116 41870
rect 45612 41410 45780 41412
rect 45612 41358 45614 41410
rect 45666 41358 45780 41410
rect 45612 41356 45780 41358
rect 45948 41858 46116 41860
rect 45948 41806 46062 41858
rect 46114 41806 46116 41858
rect 45948 41804 46116 41806
rect 45948 41410 46004 41804
rect 46060 41794 46116 41804
rect 45948 41358 45950 41410
rect 46002 41358 46004 41410
rect 45612 41346 45668 41356
rect 45948 41346 46004 41358
rect 45836 41300 45892 41310
rect 45836 41074 45892 41244
rect 45836 41022 45838 41074
rect 45890 41022 45892 41074
rect 45836 41010 45892 41022
rect 46172 40740 46228 42476
rect 46284 42466 46340 42476
rect 46396 41860 46452 41870
rect 46396 41186 46452 41804
rect 46396 41134 46398 41186
rect 46450 41134 46452 41186
rect 46396 41122 46452 41134
rect 46508 41300 46564 41310
rect 46508 40964 46564 41244
rect 45500 40684 46228 40740
rect 46396 40908 46564 40964
rect 45500 40290 45556 40684
rect 46396 40626 46452 40908
rect 46844 40740 46900 42700
rect 47180 42642 47236 42654
rect 47180 42590 47182 42642
rect 47234 42590 47236 42642
rect 47180 41300 47236 42590
rect 47180 41234 47236 41244
rect 47740 42530 47796 42542
rect 47740 42478 47742 42530
rect 47794 42478 47796 42530
rect 46844 40674 46900 40684
rect 47180 41074 47236 41086
rect 47180 41022 47182 41074
rect 47234 41022 47236 41074
rect 46396 40574 46398 40626
rect 46450 40574 46452 40626
rect 46396 40562 46452 40574
rect 46508 40628 46564 40638
rect 45500 40238 45502 40290
rect 45554 40238 45556 40290
rect 45500 40226 45556 40238
rect 46508 40290 46564 40572
rect 47180 40628 47236 41022
rect 47180 40562 47236 40572
rect 47740 40402 47796 42478
rect 48188 41858 48244 43596
rect 49308 42532 49364 42542
rect 49084 42082 49140 42094
rect 49084 42030 49086 42082
rect 49138 42030 49140 42082
rect 48748 41972 48804 41982
rect 48748 41878 48804 41916
rect 49084 41972 49140 42030
rect 48188 41806 48190 41858
rect 48242 41806 48244 41858
rect 48188 41794 48244 41806
rect 47964 40516 48020 40526
rect 47964 40422 48020 40460
rect 47740 40350 47742 40402
rect 47794 40350 47796 40402
rect 47740 40338 47796 40350
rect 48860 40404 48916 40414
rect 49084 40404 49140 41916
rect 49308 41298 49364 42476
rect 50204 42532 50260 44044
rect 50316 44034 50372 44044
rect 50428 44044 50820 44100
rect 50876 44884 50932 44894
rect 51772 44884 51828 46732
rect 51884 46722 51940 46732
rect 78204 46786 78260 46798
rect 78204 46734 78206 46786
rect 78258 46734 78260 46786
rect 78204 46452 78260 46734
rect 78204 46386 78260 46396
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 50428 42756 50484 44044
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50876 43426 50932 44828
rect 51324 44828 51828 44884
rect 51884 46004 51940 46014
rect 51324 44434 51380 44828
rect 51884 44546 51940 45948
rect 51996 45890 52052 45902
rect 51996 45838 51998 45890
rect 52050 45838 52052 45890
rect 51996 45444 52052 45838
rect 77644 45892 77700 45902
rect 77644 45798 77700 45836
rect 77420 45780 77476 45790
rect 77420 45686 77476 45724
rect 78204 45780 78260 45790
rect 78204 45686 78260 45724
rect 52668 45668 52724 45678
rect 51996 45388 52276 45444
rect 52108 45108 52164 45118
rect 52108 45014 52164 45052
rect 51884 44494 51886 44546
rect 51938 44494 51940 44546
rect 51884 44482 51940 44494
rect 51324 44382 51326 44434
rect 51378 44382 51380 44434
rect 51324 44370 51380 44382
rect 51100 44324 51156 44334
rect 51996 44324 52052 44334
rect 50988 44322 51156 44324
rect 50988 44270 51102 44322
rect 51154 44270 51156 44322
rect 50988 44268 51156 44270
rect 50988 43764 51044 44268
rect 51100 44258 51156 44268
rect 51772 44322 52052 44324
rect 51772 44270 51998 44322
rect 52050 44270 52052 44322
rect 51772 44268 52052 44270
rect 51436 44212 51492 44222
rect 51772 44212 51828 44268
rect 51996 44258 52052 44268
rect 51436 44210 51828 44212
rect 51436 44158 51438 44210
rect 51490 44158 51828 44210
rect 51436 44156 51828 44158
rect 52220 44212 52276 45388
rect 51436 43988 51492 44156
rect 52220 44146 52276 44156
rect 52668 44210 52724 45612
rect 75628 45106 75684 45118
rect 75628 45054 75630 45106
rect 75682 45054 75684 45106
rect 53340 44996 53396 45006
rect 53340 44436 53396 44940
rect 54236 44996 54292 45006
rect 54236 44902 54292 44940
rect 75404 44996 75460 45006
rect 75628 44996 75684 45054
rect 75460 44940 75684 44996
rect 77980 45108 78036 45118
rect 77980 44994 78036 45052
rect 77980 44942 77982 44994
rect 78034 44942 78036 44994
rect 75404 44902 75460 44940
rect 77980 44930 78036 44942
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 52668 44158 52670 44210
rect 52722 44158 52724 44210
rect 50988 43698 51044 43708
rect 51100 43932 51492 43988
rect 51884 44098 51940 44110
rect 51884 44046 51886 44098
rect 51938 44046 51940 44098
rect 50876 43374 50878 43426
rect 50930 43374 50932 43426
rect 50876 43362 50932 43374
rect 51100 42980 51156 43932
rect 50540 42978 51156 42980
rect 50540 42926 51102 42978
rect 51154 42926 51156 42978
rect 50540 42924 51156 42926
rect 51212 43764 51268 43774
rect 51884 43764 51940 44046
rect 51268 43708 51380 43764
rect 51212 43652 51380 43708
rect 51884 43698 51940 43708
rect 51212 42980 51268 43652
rect 51324 43540 51380 43550
rect 51324 43538 51492 43540
rect 51324 43486 51326 43538
rect 51378 43486 51492 43538
rect 51324 43484 51492 43486
rect 51324 43474 51380 43484
rect 51324 42980 51380 42990
rect 51212 42978 51380 42980
rect 51212 42926 51326 42978
rect 51378 42926 51380 42978
rect 51212 42924 51380 42926
rect 50540 42866 50596 42924
rect 51100 42914 51156 42924
rect 51324 42914 51380 42924
rect 50540 42814 50542 42866
rect 50594 42814 50596 42866
rect 50540 42802 50596 42814
rect 51436 42756 51492 43484
rect 51884 42980 51940 42990
rect 51884 42886 51940 42924
rect 50204 42466 50260 42476
rect 50316 42700 50484 42756
rect 51324 42700 51492 42756
rect 52668 42754 52724 44158
rect 52780 44434 53396 44436
rect 52780 44382 53342 44434
rect 53394 44382 53396 44434
rect 52780 44380 53396 44382
rect 52780 44210 52836 44380
rect 53340 44370 53396 44380
rect 52780 44158 52782 44210
rect 52834 44158 52836 44210
rect 52780 44146 52836 44158
rect 52892 44212 52948 44222
rect 52892 44100 52948 44156
rect 53004 44100 53060 44110
rect 52892 44098 53060 44100
rect 52892 44046 53006 44098
rect 53058 44046 53060 44098
rect 52892 44044 53060 44046
rect 53004 44034 53060 44044
rect 78204 43764 78260 43802
rect 78204 43698 78260 43708
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 52780 42980 52836 42990
rect 52780 42886 52836 42924
rect 52668 42702 52670 42754
rect 52722 42702 52724 42754
rect 50316 41972 50372 42700
rect 50652 42644 50708 42654
rect 51324 42644 51380 42700
rect 52668 42690 52724 42702
rect 51548 42644 51604 42654
rect 50652 42642 51380 42644
rect 50652 42590 50654 42642
rect 50706 42590 51380 42642
rect 50652 42588 51380 42590
rect 51436 42642 51604 42644
rect 51436 42590 51550 42642
rect 51602 42590 51604 42642
rect 51436 42588 51604 42590
rect 50652 42578 50708 42588
rect 50428 42532 50484 42542
rect 50428 42438 50484 42476
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50316 41906 50372 41916
rect 50652 41972 50708 41982
rect 50652 41878 50708 41916
rect 49308 41246 49310 41298
rect 49362 41246 49364 41298
rect 49308 41234 49364 41246
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 49532 40516 49588 40526
rect 49532 40422 49588 40460
rect 48860 40402 49140 40404
rect 48860 40350 48862 40402
rect 48914 40350 49140 40402
rect 48860 40348 49140 40350
rect 48860 40338 48916 40348
rect 46508 40238 46510 40290
rect 46562 40238 46564 40290
rect 46508 40226 46564 40238
rect 50876 40292 50932 42588
rect 51436 42082 51492 42588
rect 51548 42578 51604 42588
rect 51660 42642 51716 42654
rect 51660 42590 51662 42642
rect 51714 42590 51716 42642
rect 51660 42532 51716 42590
rect 51660 42466 51716 42476
rect 52780 42532 52836 42542
rect 53452 42532 53508 42542
rect 52780 42530 53620 42532
rect 52780 42478 52782 42530
rect 52834 42478 53454 42530
rect 53506 42478 53620 42530
rect 52780 42476 53620 42478
rect 52780 42466 52836 42476
rect 53452 42466 53508 42476
rect 51436 42030 51438 42082
rect 51490 42030 51492 42082
rect 51436 42018 51492 42030
rect 53564 41860 53620 42476
rect 77980 42420 78036 42430
rect 75628 41972 75684 41982
rect 53564 41766 53620 41804
rect 75292 41970 75684 41972
rect 75292 41918 75630 41970
rect 75682 41918 75684 41970
rect 75292 41916 75684 41918
rect 75292 41860 75348 41916
rect 75628 41906 75684 41916
rect 75292 41766 75348 41804
rect 77980 41858 78036 42364
rect 77980 41806 77982 41858
rect 78034 41806 78036 41858
rect 77980 41794 78036 41806
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 77868 41188 77924 41198
rect 77644 41076 77700 41086
rect 77644 40982 77700 41020
rect 77868 41074 77924 41132
rect 77868 41022 77870 41074
rect 77922 41022 77924 41074
rect 77868 41010 77924 41022
rect 78204 41076 78260 41086
rect 77308 40964 77364 40974
rect 75292 40628 75348 40638
rect 75348 40572 75684 40628
rect 75292 40534 75348 40572
rect 75628 40402 75684 40572
rect 77308 40514 77364 40908
rect 77308 40462 77310 40514
rect 77362 40462 77364 40514
rect 77308 40450 77364 40462
rect 75628 40350 75630 40402
rect 75682 40350 75684 40402
rect 75628 40338 75684 40350
rect 78204 40404 78260 41020
rect 78204 40338 78260 40348
rect 51660 40292 51716 40302
rect 50876 40290 51716 40292
rect 50876 40238 51662 40290
rect 51714 40238 51716 40290
rect 50876 40236 51716 40238
rect 51660 40226 51716 40236
rect 46172 40180 46228 40190
rect 45612 40178 46228 40180
rect 45612 40126 46174 40178
rect 46226 40126 46228 40178
rect 45612 40124 46228 40126
rect 45612 40068 45668 40124
rect 46172 40114 46228 40124
rect 45388 40012 45668 40068
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 44604 39554 44660 39564
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 42028 38658 42084 38668
rect 42364 38836 42420 38846
rect 40348 38612 40404 38622
rect 39844 37996 40068 38052
rect 39788 37986 39844 37996
rect 39452 37436 39732 37492
rect 39452 37266 39508 37436
rect 39452 37214 39454 37266
rect 39506 37214 39508 37266
rect 39452 37202 39508 37214
rect 39564 37266 39620 37278
rect 39564 37214 39566 37266
rect 39618 37214 39620 37266
rect 39564 36708 39620 37214
rect 39676 37266 39732 37278
rect 39676 37214 39678 37266
rect 39730 37214 39732 37266
rect 39676 37044 39732 37214
rect 39676 36978 39732 36988
rect 39564 36642 39620 36652
rect 39676 36484 39732 36494
rect 39676 36390 39732 36428
rect 40012 36482 40068 37996
rect 40348 37490 40404 38556
rect 40348 37438 40350 37490
rect 40402 37438 40404 37490
rect 40348 37426 40404 37438
rect 40012 36430 40014 36482
rect 40066 36430 40068 36482
rect 40012 36418 40068 36430
rect 40124 37266 40180 37278
rect 40124 37214 40126 37266
rect 40178 37214 40180 37266
rect 39340 36278 39396 36316
rect 39900 36258 39956 36270
rect 39900 36206 39902 36258
rect 39954 36206 39956 36258
rect 39900 35476 39956 36206
rect 39900 35410 39956 35420
rect 39340 34804 39396 34814
rect 39340 34802 39844 34804
rect 39340 34750 39342 34802
rect 39394 34750 39844 34802
rect 39340 34748 39844 34750
rect 39340 34738 39396 34748
rect 39788 34242 39844 34748
rect 39788 34190 39790 34242
rect 39842 34190 39844 34242
rect 39788 34178 39844 34190
rect 39900 34244 39956 34254
rect 39900 34130 39956 34188
rect 40124 34132 40180 37214
rect 41020 36708 41076 36718
rect 41020 36614 41076 36652
rect 40348 36482 40404 36494
rect 40348 36430 40350 36482
rect 40402 36430 40404 36482
rect 40348 36372 40404 36430
rect 40684 36484 40740 36494
rect 40684 36390 40740 36428
rect 41132 36482 41188 36494
rect 41132 36430 41134 36482
rect 41186 36430 41188 36482
rect 40348 36306 40404 36316
rect 41132 36372 41188 36430
rect 41356 36484 41412 36494
rect 41580 36484 41636 36494
rect 41412 36428 41524 36484
rect 41356 36390 41412 36428
rect 41132 36306 41188 36316
rect 39900 34078 39902 34130
rect 39954 34078 39956 34130
rect 39900 34066 39956 34078
rect 40012 34076 40180 34132
rect 40236 36258 40292 36270
rect 40236 36206 40238 36258
rect 40290 36206 40292 36258
rect 40236 34130 40292 36206
rect 41132 35476 41188 35486
rect 41188 35420 41300 35476
rect 41132 35410 41188 35420
rect 40236 34078 40238 34130
rect 40290 34078 40292 34130
rect 40012 33572 40068 34076
rect 40236 34066 40292 34078
rect 40572 34916 40628 34926
rect 40012 33506 40068 33516
rect 40124 33908 40180 33918
rect 40124 33348 40180 33852
rect 40572 33460 40628 34860
rect 40908 34916 40964 34926
rect 40908 34242 40964 34860
rect 40908 34190 40910 34242
rect 40962 34190 40964 34242
rect 40908 33908 40964 34190
rect 40908 33842 40964 33852
rect 41244 34354 41300 35420
rect 41468 35026 41524 36428
rect 41580 36390 41636 36428
rect 41804 36484 41860 36494
rect 42252 36484 42308 36494
rect 41804 36482 41972 36484
rect 41804 36430 41806 36482
rect 41858 36430 41972 36482
rect 41804 36428 41972 36430
rect 41804 36418 41860 36428
rect 41468 34974 41470 35026
rect 41522 34974 41524 35026
rect 41468 34962 41524 34974
rect 41244 34302 41246 34354
rect 41298 34302 41300 34354
rect 41244 33908 41300 34302
rect 41244 33842 41300 33852
rect 41356 34244 41412 34254
rect 41916 34244 41972 36428
rect 42252 35588 42308 36428
rect 42364 36260 42420 38780
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 78204 37826 78260 37838
rect 78204 37774 78206 37826
rect 78258 37774 78260 37826
rect 78204 37716 78260 37774
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 78204 37650 78260 37660
rect 50556 37594 50820 37604
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 42812 36596 42868 36606
rect 42812 36594 43316 36596
rect 42812 36542 42814 36594
rect 42866 36542 43316 36594
rect 42812 36540 43316 36542
rect 42812 36530 42868 36540
rect 42588 36482 42644 36494
rect 42588 36430 42590 36482
rect 42642 36430 42644 36482
rect 42588 36260 42644 36430
rect 42420 36204 42644 36260
rect 42924 36370 42980 36382
rect 42924 36318 42926 36370
rect 42978 36318 42980 36370
rect 42364 36194 42420 36204
rect 42252 34916 42308 35532
rect 42476 35698 42532 35710
rect 42476 35646 42478 35698
rect 42530 35646 42532 35698
rect 42252 34914 42420 34916
rect 42252 34862 42254 34914
rect 42306 34862 42420 34914
rect 42252 34860 42420 34862
rect 42252 34850 42308 34860
rect 42140 34244 42196 34254
rect 41916 34188 42140 34244
rect 40572 33366 40628 33404
rect 39228 33254 39284 33292
rect 39900 33292 40180 33348
rect 39788 32564 39844 32574
rect 39900 32564 39956 33292
rect 39788 32562 39956 32564
rect 39788 32510 39790 32562
rect 39842 32510 39956 32562
rect 39788 32508 39956 32510
rect 39788 32498 39844 32508
rect 40012 32452 40068 32462
rect 40012 32358 40068 32396
rect 41356 32450 41412 34188
rect 42140 34130 42196 34188
rect 42140 34078 42142 34130
rect 42194 34078 42196 34130
rect 42140 34066 42196 34078
rect 42364 34132 42420 34860
rect 42364 34038 42420 34076
rect 41804 33906 41860 33918
rect 41804 33854 41806 33906
rect 41858 33854 41860 33906
rect 41356 32398 41358 32450
rect 41410 32398 41412 32450
rect 41356 32386 41412 32398
rect 41580 33460 41636 33470
rect 41580 32564 41636 33404
rect 40348 32338 40404 32350
rect 40348 32286 40350 32338
rect 40402 32286 40404 32338
rect 39676 32004 39732 32042
rect 39676 31938 39732 31948
rect 40348 32004 40404 32286
rect 40348 31938 40404 31948
rect 39116 31780 39172 31790
rect 39564 31780 39620 31790
rect 39116 31778 39620 31780
rect 39116 31726 39118 31778
rect 39170 31726 39566 31778
rect 39618 31726 39620 31778
rect 39116 31724 39620 31726
rect 39116 31714 39172 31724
rect 39004 31556 39060 31566
rect 39004 31462 39060 31500
rect 39116 30996 39172 31006
rect 39004 30436 39060 30446
rect 38892 30380 39004 30436
rect 39004 30370 39060 30380
rect 38556 30324 38612 30334
rect 38556 30230 38612 30268
rect 38444 30158 38446 30210
rect 38498 30158 38500 30210
rect 38444 30146 38500 30158
rect 38556 29652 38612 29662
rect 38556 29558 38612 29596
rect 37884 29250 37940 29260
rect 37996 29538 38164 29540
rect 37996 29486 38110 29538
rect 38162 29486 38164 29538
rect 37996 29484 38164 29486
rect 37996 29428 38052 29484
rect 38108 29474 38164 29484
rect 37772 29204 37828 29214
rect 37548 28532 37604 28542
rect 37548 27858 37604 28476
rect 37548 27806 37550 27858
rect 37602 27806 37604 27858
rect 37548 27794 37604 27806
rect 36876 27746 37044 27748
rect 36876 27694 36878 27746
rect 36930 27694 37044 27746
rect 36876 27692 37044 27694
rect 36876 27682 36932 27692
rect 36540 27234 36596 27244
rect 36988 27074 37044 27692
rect 37100 27300 37156 27310
rect 37100 27186 37156 27244
rect 37324 27300 37380 27310
rect 37772 27300 37828 29148
rect 37884 28756 37940 28766
rect 37996 28756 38052 29372
rect 38444 29204 38500 29214
rect 38780 29204 38836 29214
rect 38332 29202 38500 29204
rect 38332 29150 38446 29202
rect 38498 29150 38500 29202
rect 38332 29148 38500 29150
rect 37884 28754 38052 28756
rect 37884 28702 37886 28754
rect 37938 28702 38052 28754
rect 37884 28700 38052 28702
rect 38220 28980 38276 28990
rect 37884 28690 37940 28700
rect 38220 28642 38276 28924
rect 38220 28590 38222 28642
rect 38274 28590 38276 28642
rect 38220 28578 38276 28590
rect 38220 27972 38276 27982
rect 38332 27972 38388 29148
rect 38444 29138 38500 29148
rect 38668 29202 38836 29204
rect 38668 29150 38782 29202
rect 38834 29150 38836 29202
rect 38668 29148 38836 29150
rect 38668 28754 38724 29148
rect 38780 29138 38836 29148
rect 38668 28702 38670 28754
rect 38722 28702 38724 28754
rect 38668 28690 38724 28702
rect 39116 28642 39172 30940
rect 39564 30884 39620 31724
rect 41020 31668 41076 31678
rect 41020 31108 41076 31612
rect 41020 31042 41076 31052
rect 41580 30996 41636 32508
rect 41804 32452 41860 33854
rect 41804 31948 41860 32396
rect 42140 33908 42196 33918
rect 41804 31892 41972 31948
rect 41916 31780 41972 31892
rect 41916 31724 42084 31780
rect 42028 31666 42084 31724
rect 42140 31778 42196 33852
rect 42476 33460 42532 35646
rect 42924 35138 42980 36318
rect 43260 35810 43316 36540
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 43260 35758 43262 35810
rect 43314 35758 43316 35810
rect 43260 35746 43316 35758
rect 45388 35588 45444 35598
rect 45388 35494 45444 35532
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 42924 35086 42926 35138
rect 42978 35086 42980 35138
rect 42924 35074 42980 35086
rect 42588 35026 42644 35038
rect 42588 34974 42590 35026
rect 42642 34974 42644 35026
rect 42588 34916 42644 34974
rect 42588 34850 42644 34860
rect 43260 34916 43316 34926
rect 42700 34244 42756 34254
rect 42700 34150 42756 34188
rect 43260 34242 43316 34860
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 43260 34190 43262 34242
rect 43314 34190 43316 34242
rect 43260 34178 43316 34190
rect 43036 34132 43092 34142
rect 43036 34038 43092 34076
rect 42476 33394 42532 33404
rect 43148 34018 43204 34030
rect 43148 33966 43150 34018
rect 43202 33966 43204 34018
rect 42140 31726 42142 31778
rect 42194 31726 42196 31778
rect 42140 31714 42196 31726
rect 42252 33124 42308 33134
rect 42028 31614 42030 31666
rect 42082 31614 42084 31666
rect 42028 31602 42084 31614
rect 41580 30902 41636 30940
rect 42140 31556 42196 31566
rect 39564 30790 39620 30828
rect 40460 30884 40516 30894
rect 39452 30436 39508 30446
rect 39452 29426 39508 30380
rect 40348 30324 40404 30334
rect 40012 30322 40404 30324
rect 40012 30270 40350 30322
rect 40402 30270 40404 30322
rect 40012 30268 40404 30270
rect 39900 30210 39956 30222
rect 39900 30158 39902 30210
rect 39954 30158 39956 30210
rect 39788 30098 39844 30110
rect 39788 30046 39790 30098
rect 39842 30046 39844 30098
rect 39452 29374 39454 29426
rect 39506 29374 39508 29426
rect 39452 29362 39508 29374
rect 39564 29986 39620 29998
rect 39564 29934 39566 29986
rect 39618 29934 39620 29986
rect 39564 29316 39620 29934
rect 39788 29988 39844 30046
rect 39564 29250 39620 29260
rect 39676 29426 39732 29438
rect 39676 29374 39678 29426
rect 39730 29374 39732 29426
rect 39452 29204 39508 29214
rect 39452 29110 39508 29148
rect 39116 28590 39118 28642
rect 39170 28590 39172 28642
rect 39116 28532 39172 28590
rect 39116 28466 39172 28476
rect 39676 28084 39732 29374
rect 39788 28980 39844 29932
rect 39900 29540 39956 30158
rect 39900 29474 39956 29484
rect 40012 29538 40068 30268
rect 40348 30258 40404 30268
rect 40460 30098 40516 30828
rect 42028 30436 42084 30446
rect 42028 30342 42084 30380
rect 41020 30324 41076 30334
rect 41020 30210 41076 30268
rect 42140 30324 42196 31500
rect 42252 30436 42308 33068
rect 43148 33012 43204 33966
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 44044 33236 44100 33246
rect 44044 33142 44100 33180
rect 45052 33236 45108 33246
rect 43820 33122 43876 33134
rect 43820 33070 43822 33122
rect 43874 33070 43876 33122
rect 43148 32956 43652 33012
rect 43484 32452 43540 32462
rect 43148 32450 43540 32452
rect 43148 32398 43486 32450
rect 43538 32398 43540 32450
rect 43148 32396 43540 32398
rect 43148 32002 43204 32396
rect 43484 32386 43540 32396
rect 43148 31950 43150 32002
rect 43202 31950 43204 32002
rect 43148 31938 43204 31950
rect 43484 31892 43540 31902
rect 43484 31798 43540 31836
rect 43596 31890 43652 32956
rect 43820 31948 43876 33070
rect 43932 33124 43988 33134
rect 43932 33030 43988 33068
rect 44156 32564 44212 32574
rect 44156 32470 44212 32508
rect 43596 31838 43598 31890
rect 43650 31838 43652 31890
rect 43596 31826 43652 31838
rect 43708 31892 43876 31948
rect 45052 32004 45108 33180
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 45052 31938 45108 31948
rect 43260 31778 43316 31790
rect 43260 31726 43262 31778
rect 43314 31726 43316 31778
rect 42364 30884 42420 30894
rect 42364 30882 42532 30884
rect 42364 30830 42366 30882
rect 42418 30830 42532 30882
rect 42364 30828 42532 30830
rect 42364 30818 42420 30828
rect 42364 30436 42420 30446
rect 42252 30434 42420 30436
rect 42252 30382 42366 30434
rect 42418 30382 42420 30434
rect 42252 30380 42420 30382
rect 42364 30370 42420 30380
rect 42196 30268 42308 30324
rect 42140 30230 42196 30268
rect 41020 30158 41022 30210
rect 41074 30158 41076 30210
rect 41020 30146 41076 30158
rect 42252 30210 42308 30268
rect 42252 30158 42254 30210
rect 42306 30158 42308 30210
rect 42252 30146 42308 30158
rect 40460 30046 40462 30098
rect 40514 30046 40516 30098
rect 40460 30034 40516 30046
rect 40684 29988 40740 29998
rect 40684 29894 40740 29932
rect 42364 29988 42420 29998
rect 42476 29988 42532 30828
rect 43260 30436 43316 31726
rect 43708 31668 43764 31892
rect 43708 31602 43764 31612
rect 44828 31778 44884 31790
rect 44828 31726 44830 31778
rect 44882 31726 44884 31778
rect 44828 31668 44884 31726
rect 44492 30884 44548 30894
rect 44828 30884 44884 31612
rect 45388 31556 45444 31566
rect 45388 31462 45444 31500
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 44492 30882 44884 30884
rect 44492 30830 44494 30882
rect 44546 30830 44884 30882
rect 44492 30828 44884 30830
rect 44492 30818 44548 30828
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 43260 30370 43316 30380
rect 42364 29986 42532 29988
rect 42364 29934 42366 29986
rect 42418 29934 42532 29986
rect 42364 29932 42532 29934
rect 78204 30322 78260 30334
rect 78204 30270 78206 30322
rect 78258 30270 78260 30322
rect 42364 29922 42420 29932
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 78204 29764 78260 30270
rect 78204 29698 78260 29708
rect 40012 29486 40014 29538
rect 40066 29486 40068 29538
rect 40012 29474 40068 29486
rect 41020 29540 41076 29550
rect 39788 28914 39844 28924
rect 39900 29314 39956 29326
rect 39900 29262 39902 29314
rect 39954 29262 39956 29314
rect 39788 28756 39844 28766
rect 39900 28756 39956 29262
rect 39788 28754 39956 28756
rect 39788 28702 39790 28754
rect 39842 28702 39956 28754
rect 39788 28700 39956 28702
rect 40348 28980 40404 28990
rect 39788 28690 39844 28700
rect 39676 28018 39732 28028
rect 38220 27970 38388 27972
rect 38220 27918 38222 27970
rect 38274 27918 38388 27970
rect 38220 27916 38388 27918
rect 38220 27906 38276 27916
rect 40348 27746 40404 28924
rect 41020 28756 41076 29484
rect 78204 29538 78260 29550
rect 78204 29486 78206 29538
rect 78258 29486 78260 29538
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 78204 28980 78260 29486
rect 78204 28914 78260 28924
rect 40908 28084 40964 28094
rect 40908 27990 40964 28028
rect 41020 27970 41076 28700
rect 41916 28756 41972 28766
rect 41916 28662 41972 28700
rect 78204 28418 78260 28430
rect 78204 28366 78206 28418
rect 78258 28366 78260 28418
rect 78204 28308 78260 28366
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 78204 28242 78260 28252
rect 50556 28186 50820 28196
rect 41020 27918 41022 27970
rect 41074 27918 41076 27970
rect 41020 27906 41076 27918
rect 40348 27694 40350 27746
rect 40402 27694 40404 27746
rect 40348 27682 40404 27694
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 37324 27298 37828 27300
rect 37324 27246 37326 27298
rect 37378 27246 37828 27298
rect 37324 27244 37828 27246
rect 37324 27234 37380 27244
rect 37100 27134 37102 27186
rect 37154 27134 37156 27186
rect 37100 27122 37156 27134
rect 78204 27186 78260 27198
rect 78204 27134 78206 27186
rect 78258 27134 78260 27186
rect 36988 27022 36990 27074
rect 37042 27022 37044 27074
rect 36988 27010 37044 27022
rect 78204 26964 78260 27134
rect 78204 26898 78260 26908
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 78204 20244 78260 20282
rect 36316 20132 36484 20188
rect 78204 20178 78260 20188
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 28252 4228 28308 4238
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 28252 800 28308 4172
rect 36428 4228 36484 20132
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 78204 19346 78260 19358
rect 78204 19294 78206 19346
rect 78258 19294 78260 19346
rect 78204 18900 78260 19294
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 78204 18834 78260 18844
rect 50556 18778 50820 18788
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 78204 17444 78260 17454
rect 78204 17442 78372 17444
rect 78204 17390 78206 17442
rect 78258 17390 78372 17442
rect 78204 17388 78372 17390
rect 78204 17378 78260 17388
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 78204 16994 78260 17006
rect 78204 16942 78206 16994
rect 78258 16942 78260 16994
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 78204 16212 78260 16942
rect 78316 16884 78372 17388
rect 78428 16884 78484 16894
rect 78316 16828 78428 16884
rect 78428 16818 78484 16828
rect 78204 16146 78260 16156
rect 78204 15874 78260 15886
rect 78204 15822 78206 15874
rect 78258 15822 78260 15874
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 78204 15540 78260 15822
rect 78204 15474 78260 15484
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 36428 4162 36484 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 35196 3332 35252 3342
rect 38556 3332 38612 3342
rect 48636 3332 48692 3342
rect 49980 3332 50036 3342
rect 59388 3332 59444 3342
rect 62748 3332 62804 3342
rect 63420 3332 63476 3342
rect 67452 3332 67508 3342
rect 34972 3330 35252 3332
rect 34972 3278 35198 3330
rect 35250 3278 35252 3330
rect 34972 3276 35252 3278
rect 34972 800 35028 3276
rect 35196 3266 35252 3276
rect 38332 3330 38612 3332
rect 38332 3278 38558 3330
rect 38610 3278 38612 3330
rect 38332 3276 38612 3278
rect 38332 800 38388 3276
rect 38556 3266 38612 3276
rect 48412 3330 48692 3332
rect 48412 3278 48638 3330
rect 48690 3278 48692 3330
rect 48412 3276 48692 3278
rect 48412 800 48468 3276
rect 48636 3266 48692 3276
rect 49756 3330 50036 3332
rect 49756 3278 49982 3330
rect 50034 3278 50036 3330
rect 49756 3276 50036 3278
rect 49756 800 49812 3276
rect 49980 3266 50036 3276
rect 59164 3330 59444 3332
rect 59164 3278 59390 3330
rect 59442 3278 59444 3330
rect 59164 3276 59444 3278
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 59164 800 59220 3276
rect 59388 3266 59444 3276
rect 62524 3330 62804 3332
rect 62524 3278 62750 3330
rect 62802 3278 62804 3330
rect 62524 3276 62804 3278
rect 62524 800 62580 3276
rect 62748 3266 62804 3276
rect 63196 3330 63476 3332
rect 63196 3278 63422 3330
rect 63474 3278 63476 3330
rect 63196 3276 63476 3278
rect 63196 800 63252 3276
rect 63420 3266 63476 3276
rect 67228 3330 67508 3332
rect 67228 3278 67454 3330
rect 67506 3278 67508 3330
rect 67228 3276 67508 3278
rect 67228 800 67284 3276
rect 67452 3266 67508 3276
rect 28224 0 28336 800
rect 34944 0 35056 800
rect 38304 0 38416 800
rect 48384 0 48496 800
rect 49728 0 49840 800
rect 59136 0 59248 800
rect 62496 0 62608 800
rect 63168 0 63280 800
rect 67200 0 67312 800
<< via2 >>
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 78204 64594 78260 64596
rect 78204 64542 78206 64594
rect 78206 64542 78258 64594
rect 78258 64542 78260 64594
rect 78204 64540 78260 64542
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 78204 60562 78260 60564
rect 78204 60510 78206 60562
rect 78206 60510 78258 60562
rect 78258 60510 78260 60562
rect 78204 60508 78260 60510
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 78204 59890 78260 59892
rect 78204 59838 78206 59890
rect 78206 59838 78258 59890
rect 78258 59838 78260 59890
rect 78204 59836 78260 59838
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 78204 57820 78260 57876
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 47852 49138 47908 49140
rect 47852 49086 47854 49138
rect 47854 49086 47906 49138
rect 47906 49086 47908 49138
rect 47852 49084 47908 49086
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 29148 47180 29204 47236
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 30492 47234 30548 47236
rect 30492 47182 30494 47234
rect 30494 47182 30546 47234
rect 30546 47182 30548 47234
rect 30492 47180 30548 47182
rect 30380 47068 30436 47124
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 28476 45836 28532 45892
rect 29260 45890 29316 45892
rect 29260 45838 29262 45890
rect 29262 45838 29314 45890
rect 29314 45838 29316 45890
rect 29260 45836 29316 45838
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 29932 45276 29988 45332
rect 31276 46562 31332 46564
rect 31276 46510 31278 46562
rect 31278 46510 31330 46562
rect 31330 46510 31332 46562
rect 31276 46508 31332 46510
rect 31612 45276 31668 45332
rect 31948 46508 32004 46564
rect 32396 45836 32452 45892
rect 32172 45612 32228 45668
rect 30828 44828 30884 44884
rect 29932 43260 29988 43316
rect 30716 43314 30772 43316
rect 30716 43262 30718 43314
rect 30718 43262 30770 43314
rect 30770 43262 30772 43314
rect 30716 43260 30772 43262
rect 31724 44882 31780 44884
rect 31724 44830 31726 44882
rect 31726 44830 31778 44882
rect 31778 44830 31780 44882
rect 31724 44828 31780 44830
rect 30940 43596 30996 43652
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 28028 41804 28084 41860
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 32060 42700 32116 42756
rect 32508 42700 32564 42756
rect 29260 41804 29316 41860
rect 29708 41804 29764 41860
rect 28700 41356 28756 41412
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 30604 41410 30660 41412
rect 30604 41358 30606 41410
rect 30606 41358 30658 41410
rect 30658 41358 30660 41410
rect 30604 41356 30660 41358
rect 30828 41916 30884 41972
rect 31724 41970 31780 41972
rect 31724 41918 31726 41970
rect 31726 41918 31778 41970
rect 31778 41918 31780 41970
rect 31724 41916 31780 41918
rect 32396 41970 32452 41972
rect 32396 41918 32398 41970
rect 32398 41918 32450 41970
rect 32450 41918 32452 41970
rect 32396 41916 32452 41918
rect 31500 41746 31556 41748
rect 31500 41694 31502 41746
rect 31502 41694 31554 41746
rect 31554 41694 31556 41746
rect 31500 41692 31556 41694
rect 32060 41746 32116 41748
rect 32060 41694 32062 41746
rect 32062 41694 32114 41746
rect 32114 41694 32116 41746
rect 32060 41692 32116 41694
rect 31164 41356 31220 41412
rect 30380 40236 30436 40292
rect 30716 40236 30772 40292
rect 31164 40348 31220 40404
rect 31500 40012 31556 40068
rect 32172 41356 32228 41412
rect 34636 47068 34692 47124
rect 33068 46508 33124 46564
rect 33292 45890 33348 45892
rect 33292 45838 33294 45890
rect 33294 45838 33346 45890
rect 33346 45838 33348 45890
rect 33292 45836 33348 45838
rect 33180 45612 33236 45668
rect 33628 45276 33684 45332
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 34076 45666 34132 45668
rect 34076 45614 34078 45666
rect 34078 45614 34130 45666
rect 34130 45614 34132 45666
rect 34076 45612 34132 45614
rect 34412 45276 34468 45332
rect 34300 45218 34356 45220
rect 34300 45166 34302 45218
rect 34302 45166 34354 45218
rect 34354 45166 34356 45218
rect 34300 45164 34356 45166
rect 33852 44828 33908 44884
rect 33964 45052 34020 45108
rect 34300 43650 34356 43652
rect 34300 43598 34302 43650
rect 34302 43598 34354 43650
rect 34354 43598 34356 43650
rect 34300 43596 34356 43598
rect 33404 42700 33460 42756
rect 32956 41804 33012 41860
rect 32060 40348 32116 40404
rect 32060 40012 32116 40068
rect 32396 39842 32452 39844
rect 32396 39790 32398 39842
rect 32398 39790 32450 39842
rect 32450 39790 32452 39842
rect 32396 39788 32452 39790
rect 31836 39452 31892 39508
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 30156 37996 30212 38052
rect 29148 36988 29204 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 28140 31836 28196 31892
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 32508 39676 32564 39732
rect 32620 39452 32676 39508
rect 32956 40012 33012 40068
rect 32956 39842 33012 39844
rect 32956 39790 32958 39842
rect 32958 39790 33010 39842
rect 33010 39790 33012 39842
rect 32956 39788 33012 39790
rect 34636 45164 34692 45220
rect 35084 45612 35140 45668
rect 35420 45836 35476 45892
rect 35308 45276 35364 45332
rect 34748 45106 34804 45108
rect 34748 45054 34750 45106
rect 34750 45054 34802 45106
rect 34802 45054 34804 45106
rect 34748 45052 34804 45054
rect 34972 45052 35028 45108
rect 34748 44828 34804 44884
rect 35644 45724 35700 45780
rect 35532 45164 35588 45220
rect 38556 46620 38612 46676
rect 36988 45890 37044 45892
rect 36988 45838 36990 45890
rect 36990 45838 37042 45890
rect 37042 45838 37044 45890
rect 36988 45836 37044 45838
rect 36428 45724 36484 45780
rect 35868 45164 35924 45220
rect 36316 45218 36372 45220
rect 36316 45166 36318 45218
rect 36318 45166 36370 45218
rect 36370 45166 36372 45218
rect 36316 45164 36372 45166
rect 36428 45106 36484 45108
rect 36428 45054 36430 45106
rect 36430 45054 36482 45106
rect 36482 45054 36484 45106
rect 36428 45052 36484 45054
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35532 44546 35588 44548
rect 35532 44494 35534 44546
rect 35534 44494 35586 44546
rect 35586 44494 35588 44546
rect 35532 44492 35588 44494
rect 37212 44492 37268 44548
rect 34860 43596 34916 43652
rect 36316 43484 36372 43540
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 33852 42530 33908 42532
rect 33852 42478 33854 42530
rect 33854 42478 33906 42530
rect 33906 42478 33908 42530
rect 33852 42476 33908 42478
rect 33740 41916 33796 41972
rect 34972 42028 35028 42084
rect 33516 41858 33572 41860
rect 33516 41806 33518 41858
rect 33518 41806 33570 41858
rect 33570 41806 33572 41858
rect 33516 41804 33572 41806
rect 34636 40514 34692 40516
rect 34636 40462 34638 40514
rect 34638 40462 34690 40514
rect 34690 40462 34692 40514
rect 34636 40460 34692 40462
rect 34300 40236 34356 40292
rect 33180 39506 33236 39508
rect 33180 39454 33182 39506
rect 33182 39454 33234 39506
rect 33234 39454 33236 39506
rect 33180 39452 33236 39454
rect 37212 42866 37268 42868
rect 37212 42814 37214 42866
rect 37214 42814 37266 42866
rect 37266 42814 37268 42866
rect 37212 42812 37268 42814
rect 36428 42754 36484 42756
rect 36428 42702 36430 42754
rect 36430 42702 36482 42754
rect 36482 42702 36484 42754
rect 36428 42700 36484 42702
rect 37436 42754 37492 42756
rect 37436 42702 37438 42754
rect 37438 42702 37490 42754
rect 37490 42702 37492 42754
rect 37436 42700 37492 42702
rect 37660 42028 37716 42084
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35756 41020 35812 41076
rect 37436 41020 37492 41076
rect 42028 46620 42084 46676
rect 39564 45276 39620 45332
rect 37884 44268 37940 44324
rect 38668 44882 38724 44884
rect 38668 44830 38670 44882
rect 38670 44830 38722 44882
rect 38722 44830 38724 44882
rect 38668 44828 38724 44830
rect 39004 44604 39060 44660
rect 40348 45276 40404 45332
rect 39564 44604 39620 44660
rect 39788 44828 39844 44884
rect 39228 44492 39284 44548
rect 39564 44322 39620 44324
rect 39564 44270 39566 44322
rect 39566 44270 39618 44322
rect 39618 44270 39620 44322
rect 39564 44268 39620 44270
rect 38444 43820 38500 43876
rect 38444 43596 38500 43652
rect 38668 43484 38724 43540
rect 38108 42700 38164 42756
rect 38220 42812 38276 42868
rect 38332 41916 38388 41972
rect 38556 42140 38612 42196
rect 38444 41804 38500 41860
rect 38668 41410 38724 41412
rect 38668 41358 38670 41410
rect 38670 41358 38722 41410
rect 38722 41358 38724 41410
rect 38668 41356 38724 41358
rect 38892 42476 38948 42532
rect 39116 42028 39172 42084
rect 39452 43596 39508 43652
rect 41132 45276 41188 45332
rect 43036 46562 43092 46564
rect 43036 46510 43038 46562
rect 43038 46510 43090 46562
rect 43090 46510 43092 46562
rect 43036 46508 43092 46510
rect 39900 43484 39956 43540
rect 39564 43036 39620 43092
rect 39452 41356 39508 41412
rect 38780 41132 38836 41188
rect 39564 41132 39620 41188
rect 37772 40572 37828 40628
rect 39228 40572 39284 40628
rect 35756 40460 35812 40516
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 37100 40514 37156 40516
rect 37100 40462 37102 40514
rect 37102 40462 37154 40514
rect 37154 40462 37156 40514
rect 37100 40460 37156 40462
rect 37884 40402 37940 40404
rect 37884 40350 37886 40402
rect 37886 40350 37938 40402
rect 37938 40350 37940 40402
rect 37884 40348 37940 40350
rect 39004 40012 39060 40068
rect 35532 38668 35588 38724
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35084 37996 35140 38052
rect 34300 37884 34356 37940
rect 33628 36988 33684 37044
rect 35420 37938 35476 37940
rect 35420 37886 35422 37938
rect 35422 37886 35474 37938
rect 35474 37886 35476 37938
rect 35420 37884 35476 37886
rect 34748 36988 34804 37044
rect 31500 36204 31556 36260
rect 29932 34802 29988 34804
rect 29932 34750 29934 34802
rect 29934 34750 29986 34802
rect 29986 34750 29988 34802
rect 29932 34748 29988 34750
rect 31388 34748 31444 34804
rect 32172 36258 32228 36260
rect 32172 36206 32174 36258
rect 32174 36206 32226 36258
rect 32226 36206 32228 36258
rect 32172 36204 32228 36206
rect 31276 33404 31332 33460
rect 31724 33906 31780 33908
rect 31724 33854 31726 33906
rect 31726 33854 31778 33906
rect 31778 33854 31780 33906
rect 31724 33852 31780 33854
rect 30940 33180 30996 33236
rect 29148 31836 29204 31892
rect 28812 31500 28868 31556
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 30604 31554 30660 31556
rect 30604 31502 30606 31554
rect 30606 31502 30658 31554
rect 30658 31502 30660 31554
rect 30604 31500 30660 31502
rect 31612 33234 31668 33236
rect 31612 33182 31614 33234
rect 31614 33182 31666 33234
rect 31666 33182 31668 33234
rect 31612 33180 31668 33182
rect 32172 33346 32228 33348
rect 32172 33294 32174 33346
rect 32174 33294 32226 33346
rect 32226 33294 32228 33346
rect 32172 33292 32228 33294
rect 33852 33906 33908 33908
rect 33852 33854 33854 33906
rect 33854 33854 33906 33906
rect 33906 33854 33908 33906
rect 33852 33852 33908 33854
rect 33404 33404 33460 33460
rect 32396 33292 32452 33348
rect 31948 32956 32004 33012
rect 31500 31890 31556 31892
rect 31500 31838 31502 31890
rect 31502 31838 31554 31890
rect 31554 31838 31556 31890
rect 31500 31836 31556 31838
rect 32172 32844 32228 32900
rect 32172 31836 32228 31892
rect 32284 31164 32340 31220
rect 32396 32284 32452 32340
rect 33516 32284 33572 32340
rect 34076 32956 34132 33012
rect 33964 32844 34020 32900
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35532 36652 35588 36708
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36988 38722 37044 38724
rect 36988 38670 36990 38722
rect 36990 38670 37042 38722
rect 37042 38670 37044 38722
rect 36988 38668 37044 38670
rect 35756 38050 35812 38052
rect 35756 37998 35758 38050
rect 35758 37998 35810 38050
rect 35810 37998 35812 38050
rect 35756 37996 35812 37998
rect 35980 38050 36036 38052
rect 35980 37998 35982 38050
rect 35982 37998 36034 38050
rect 36034 37998 36036 38050
rect 35980 37996 36036 37998
rect 36428 36876 36484 36932
rect 35644 34300 35700 34356
rect 36204 34300 36260 34356
rect 35084 33852 35140 33908
rect 34748 33458 34804 33460
rect 34748 33406 34750 33458
rect 34750 33406 34802 33458
rect 34802 33406 34804 33458
rect 34748 33404 34804 33406
rect 34972 33346 35028 33348
rect 34972 33294 34974 33346
rect 34974 33294 35026 33346
rect 35026 33294 35028 33346
rect 34972 33292 35028 33294
rect 34300 31218 34356 31220
rect 34300 31166 34302 31218
rect 34302 31166 34354 31218
rect 34354 31166 34356 31218
rect 34300 31164 34356 31166
rect 32508 30828 32564 30884
rect 33628 30882 33684 30884
rect 33628 30830 33630 30882
rect 33630 30830 33682 30882
rect 33682 30830 33684 30882
rect 33628 30828 33684 30830
rect 30492 30268 30548 30324
rect 31388 30268 31444 30324
rect 30156 29148 30212 29204
rect 31276 29202 31332 29204
rect 31276 29150 31278 29202
rect 31278 29150 31330 29202
rect 31330 29150 31332 29202
rect 31276 29148 31332 29150
rect 29372 28642 29428 28644
rect 29372 28590 29374 28642
rect 29374 28590 29426 28642
rect 29426 28590 29428 28642
rect 29372 28588 29428 28590
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 32172 29148 32228 29204
rect 33516 29426 33572 29428
rect 33516 29374 33518 29426
rect 33518 29374 33570 29426
rect 33570 29374 33572 29426
rect 33516 29372 33572 29374
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35980 33122 36036 33124
rect 35980 33070 35982 33122
rect 35982 33070 36034 33122
rect 36034 33070 36036 33122
rect 35980 33068 36036 33070
rect 35980 31612 36036 31668
rect 36092 31500 36148 31556
rect 36316 31106 36372 31108
rect 36316 31054 36318 31106
rect 36318 31054 36370 31106
rect 36370 31054 36372 31106
rect 36316 31052 36372 31054
rect 36988 36706 37044 36708
rect 36988 36654 36990 36706
rect 36990 36654 37042 36706
rect 37042 36654 37044 36706
rect 36988 36652 37044 36654
rect 37324 36876 37380 36932
rect 39228 38108 39284 38164
rect 38556 37996 38612 38052
rect 37996 36988 38052 37044
rect 38220 36876 38276 36932
rect 39116 36764 39172 36820
rect 37660 36540 37716 36596
rect 38892 36594 38948 36596
rect 38892 36542 38894 36594
rect 38894 36542 38946 36594
rect 38946 36542 38948 36594
rect 38892 36540 38948 36542
rect 37324 36370 37380 36372
rect 37324 36318 37326 36370
rect 37326 36318 37378 36370
rect 37378 36318 37380 36370
rect 37324 36316 37380 36318
rect 37100 34354 37156 34356
rect 37100 34302 37102 34354
rect 37102 34302 37154 34354
rect 37154 34302 37156 34354
rect 37100 34300 37156 34302
rect 37436 34242 37492 34244
rect 37436 34190 37438 34242
rect 37438 34190 37490 34242
rect 37490 34190 37492 34242
rect 37436 34188 37492 34190
rect 36764 30994 36820 30996
rect 36764 30942 36766 30994
rect 36766 30942 36818 30994
rect 36818 30942 36820 30994
rect 36764 30940 36820 30942
rect 35196 29426 35252 29428
rect 35196 29374 35198 29426
rect 35198 29374 35250 29426
rect 35250 29374 35252 29426
rect 35196 29372 35252 29374
rect 33740 29202 33796 29204
rect 33740 29150 33742 29202
rect 33742 29150 33794 29202
rect 33794 29150 33796 29202
rect 33740 29148 33796 29150
rect 33852 28812 33908 28868
rect 32620 28642 32676 28644
rect 32620 28590 32622 28642
rect 32622 28590 32674 28642
rect 32674 28590 32676 28642
rect 32620 28588 32676 28590
rect 33964 28588 34020 28644
rect 35420 29202 35476 29204
rect 35420 29150 35422 29202
rect 35422 29150 35474 29202
rect 35474 29150 35476 29202
rect 35420 29148 35476 29150
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 36204 30380 36260 30436
rect 36204 29596 36260 29652
rect 35980 28812 36036 28868
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 36988 30380 37044 30436
rect 37100 31666 37156 31668
rect 37100 31614 37102 31666
rect 37102 31614 37154 31666
rect 37154 31614 37156 31666
rect 37100 31612 37156 31614
rect 37212 31164 37268 31220
rect 37548 33122 37604 33124
rect 37548 33070 37550 33122
rect 37550 33070 37602 33122
rect 37602 33070 37604 33122
rect 37548 33068 37604 33070
rect 37100 29650 37156 29652
rect 37100 29598 37102 29650
rect 37102 29598 37154 29650
rect 37154 29598 37156 29650
rect 37100 29596 37156 29598
rect 37548 30268 37604 30324
rect 38668 34914 38724 34916
rect 38668 34862 38670 34914
rect 38670 34862 38722 34914
rect 38722 34862 38724 34914
rect 38668 34860 38724 34862
rect 38892 34188 38948 34244
rect 38332 33292 38388 33348
rect 38556 31948 38612 32004
rect 37772 29596 37828 29652
rect 36652 29426 36708 29428
rect 36652 29374 36654 29426
rect 36654 29374 36706 29426
rect 36706 29374 36708 29426
rect 36652 29372 36708 29374
rect 36428 29314 36484 29316
rect 36428 29262 36430 29314
rect 36430 29262 36482 29314
rect 36482 29262 36484 29314
rect 36428 29260 36484 29262
rect 36540 29148 36596 29204
rect 38444 31500 38500 31556
rect 39564 38162 39620 38164
rect 39564 38110 39566 38162
rect 39566 38110 39618 38162
rect 39618 38110 39620 38162
rect 39564 38108 39620 38110
rect 40348 43036 40404 43092
rect 43372 44940 43428 44996
rect 42140 44210 42196 44212
rect 42140 44158 42142 44210
rect 42142 44158 42194 44210
rect 42194 44158 42196 44210
rect 42140 44156 42196 44158
rect 47628 48466 47684 48468
rect 47628 48414 47630 48466
rect 47630 48414 47682 48466
rect 47682 48414 47684 48466
rect 47628 48412 47684 48414
rect 47740 48354 47796 48356
rect 47740 48302 47742 48354
rect 47742 48302 47794 48354
rect 47794 48302 47796 48354
rect 47740 48300 47796 48302
rect 46284 47964 46340 48020
rect 46284 47180 46340 47236
rect 45836 47068 45892 47124
rect 46844 47292 46900 47348
rect 46620 47234 46676 47236
rect 46620 47182 46622 47234
rect 46622 47182 46674 47234
rect 46674 47182 46676 47234
rect 46620 47180 46676 47182
rect 46732 47068 46788 47124
rect 45500 46620 45556 46676
rect 45276 45164 45332 45220
rect 44940 44098 44996 44100
rect 44940 44046 44942 44098
rect 44942 44046 44994 44098
rect 44994 44046 44996 44098
rect 44940 44044 44996 44046
rect 40796 41970 40852 41972
rect 40796 41918 40798 41970
rect 40798 41918 40850 41970
rect 40850 41918 40852 41970
rect 40796 41916 40852 41918
rect 41132 41970 41188 41972
rect 41132 41918 41134 41970
rect 41134 41918 41186 41970
rect 41186 41918 41188 41970
rect 41132 41916 41188 41918
rect 39900 41244 39956 41300
rect 41244 41298 41300 41300
rect 41244 41246 41246 41298
rect 41246 41246 41298 41298
rect 41298 41246 41300 41298
rect 41244 41244 41300 41246
rect 41020 40460 41076 40516
rect 41468 41132 41524 41188
rect 45388 44210 45444 44212
rect 45388 44158 45390 44210
rect 45390 44158 45442 44210
rect 45442 44158 45444 44210
rect 45388 44156 45444 44158
rect 46396 46674 46452 46676
rect 46396 46622 46398 46674
rect 46398 46622 46450 46674
rect 46450 46622 46452 46674
rect 46396 46620 46452 46622
rect 46508 46562 46564 46564
rect 46508 46510 46510 46562
rect 46510 46510 46562 46562
rect 46562 46510 46564 46562
rect 46508 46508 46564 46510
rect 47180 46114 47236 46116
rect 47180 46062 47182 46114
rect 47182 46062 47234 46114
rect 47234 46062 47236 46114
rect 47180 46060 47236 46062
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 78204 49756 78260 49812
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 49532 49084 49588 49140
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 48748 48466 48804 48468
rect 48748 48414 48750 48466
rect 48750 48414 48802 48466
rect 48802 48414 48804 48466
rect 48748 48412 48804 48414
rect 47852 47964 47908 48020
rect 47740 47346 47796 47348
rect 47740 47294 47742 47346
rect 47742 47294 47794 47346
rect 47794 47294 47796 47346
rect 47740 47292 47796 47294
rect 47516 47068 47572 47124
rect 47628 46956 47684 47012
rect 47404 46620 47460 46676
rect 47740 46674 47796 46676
rect 47740 46622 47742 46674
rect 47742 46622 47794 46674
rect 47794 46622 47796 46674
rect 47740 46620 47796 46622
rect 47628 46508 47684 46564
rect 47516 46396 47572 46452
rect 48188 47404 48244 47460
rect 48300 47180 48356 47236
rect 48300 46786 48356 46788
rect 48300 46734 48302 46786
rect 48302 46734 48354 46786
rect 48354 46734 48356 46786
rect 48300 46732 48356 46734
rect 49756 48300 49812 48356
rect 49084 48242 49140 48244
rect 49084 48190 49086 48242
rect 49086 48190 49138 48242
rect 49138 48190 49140 48242
rect 49084 48188 49140 48190
rect 49532 48130 49588 48132
rect 49532 48078 49534 48130
rect 49534 48078 49586 48130
rect 49586 48078 49588 48130
rect 49532 48076 49588 48078
rect 48748 47516 48804 47572
rect 48636 47234 48692 47236
rect 48636 47182 48638 47234
rect 48638 47182 48690 47234
rect 48690 47182 48692 47234
rect 48636 47180 48692 47182
rect 48524 46620 48580 46676
rect 46060 45218 46116 45220
rect 46060 45166 46062 45218
rect 46062 45166 46114 45218
rect 46114 45166 46116 45218
rect 46060 45164 46116 45166
rect 45836 45106 45892 45108
rect 45836 45054 45838 45106
rect 45838 45054 45890 45106
rect 45890 45054 45892 45106
rect 45836 45052 45892 45054
rect 45948 44994 46004 44996
rect 45948 44942 45950 44994
rect 45950 44942 46002 44994
rect 46002 44942 46004 44994
rect 45948 44940 46004 44942
rect 48748 46674 48804 46676
rect 48748 46622 48750 46674
rect 48750 46622 48802 46674
rect 48802 46622 48804 46674
rect 48748 46620 48804 46622
rect 48636 46508 48692 46564
rect 48860 46450 48916 46452
rect 48860 46398 48862 46450
rect 48862 46398 48914 46450
rect 48914 46398 48916 46450
rect 48860 46396 48916 46398
rect 49196 47458 49252 47460
rect 49196 47406 49198 47458
rect 49198 47406 49250 47458
rect 49250 47406 49252 47458
rect 49196 47404 49252 47406
rect 49420 47516 49476 47572
rect 49980 48188 50036 48244
rect 49420 46844 49476 46900
rect 49084 46786 49140 46788
rect 49084 46734 49086 46786
rect 49086 46734 49138 46786
rect 49138 46734 49140 46786
rect 49084 46732 49140 46734
rect 46956 45500 47012 45556
rect 48636 45724 48692 45780
rect 48076 45666 48132 45668
rect 48076 45614 48078 45666
rect 48078 45614 48130 45666
rect 48130 45614 48132 45666
rect 48076 45612 48132 45614
rect 49420 46172 49476 46228
rect 50540 48130 50596 48132
rect 50540 48078 50542 48130
rect 50542 48078 50594 48130
rect 50594 48078 50596 48130
rect 50540 48076 50596 48078
rect 50540 47628 50596 47684
rect 51100 47628 51156 47684
rect 50204 46956 50260 47012
rect 49980 46620 50036 46676
rect 49868 46396 49924 46452
rect 49756 46060 49812 46116
rect 47964 45276 48020 45332
rect 47068 45106 47124 45108
rect 47068 45054 47070 45106
rect 47070 45054 47122 45106
rect 47122 45054 47124 45106
rect 47068 45052 47124 45054
rect 49420 45612 49476 45668
rect 47852 44994 47908 44996
rect 47852 44942 47854 44994
rect 47854 44942 47906 44994
rect 47906 44942 47908 44994
rect 47852 44940 47908 44942
rect 48860 45330 48916 45332
rect 48860 45278 48862 45330
rect 48862 45278 48914 45330
rect 48914 45278 48916 45330
rect 48860 45276 48916 45278
rect 49868 45500 49924 45556
rect 50316 46786 50372 46788
rect 50316 46734 50318 46786
rect 50318 46734 50370 46786
rect 50370 46734 50372 46786
rect 50316 46732 50372 46734
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50876 46674 50932 46676
rect 50876 46622 50878 46674
rect 50878 46622 50930 46674
rect 50930 46622 50932 46674
rect 50876 46620 50932 46622
rect 50876 45948 50932 46004
rect 51100 46898 51156 46900
rect 51100 46846 51102 46898
rect 51102 46846 51154 46898
rect 51154 46846 51156 46898
rect 51100 46844 51156 46846
rect 50988 46172 51044 46228
rect 50652 45890 50708 45892
rect 50652 45838 50654 45890
rect 50654 45838 50706 45890
rect 50706 45838 50708 45890
rect 50652 45836 50708 45838
rect 50316 45724 50372 45780
rect 48636 44940 48692 44996
rect 49868 44546 49924 44548
rect 49868 44494 49870 44546
rect 49870 44494 49922 44546
rect 49922 44494 49924 44546
rect 49868 44492 49924 44494
rect 43036 41244 43092 41300
rect 41692 41020 41748 41076
rect 42252 41132 42308 41188
rect 42028 40796 42084 40852
rect 41132 40012 41188 40068
rect 42028 39564 42084 39620
rect 41132 38780 41188 38836
rect 42812 41186 42868 41188
rect 42812 41134 42814 41186
rect 42814 41134 42866 41186
rect 42866 41134 42868 41186
rect 42812 41132 42868 41134
rect 44156 41244 44212 41300
rect 43484 41186 43540 41188
rect 43484 41134 43486 41186
rect 43486 41134 43538 41186
rect 43538 41134 43540 41186
rect 43484 41132 43540 41134
rect 43372 40908 43428 40964
rect 42700 40796 42756 40852
rect 43932 40962 43988 40964
rect 43932 40910 43934 40962
rect 43934 40910 43986 40962
rect 43986 40910 43988 40962
rect 43932 40908 43988 40910
rect 42924 39564 42980 39620
rect 43260 39618 43316 39620
rect 43260 39566 43262 39618
rect 43262 39566 43314 39618
rect 43314 39566 43316 39618
rect 43260 39564 43316 39566
rect 44940 41970 44996 41972
rect 44940 41918 44942 41970
rect 44942 41918 44994 41970
rect 44994 41918 44996 41970
rect 44940 41916 44996 41918
rect 45724 44044 45780 44100
rect 45276 41804 45332 41860
rect 45500 42924 45556 42980
rect 45612 41916 45668 41972
rect 49756 43708 49812 43764
rect 51772 47346 51828 47348
rect 51772 47294 51774 47346
rect 51774 47294 51826 47346
rect 51826 47294 51828 47346
rect 51772 47292 51828 47294
rect 51436 46844 51492 46900
rect 52668 47346 52724 47348
rect 52668 47294 52670 47346
rect 52670 47294 52722 47346
rect 52722 47294 52724 47346
rect 52668 47292 52724 47294
rect 52892 47292 52948 47348
rect 53340 47346 53396 47348
rect 53340 47294 53342 47346
rect 53342 47294 53394 47346
rect 53394 47294 53396 47346
rect 53340 47292 53396 47294
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 53676 47292 53732 47348
rect 77980 47740 78036 47796
rect 75404 47292 75460 47348
rect 77868 47628 77924 47684
rect 77644 47068 77700 47124
rect 78204 47068 78260 47124
rect 51884 46732 51940 46788
rect 51436 45778 51492 45780
rect 51436 45726 51438 45778
rect 51438 45726 51490 45778
rect 51490 45726 51492 45778
rect 51436 45724 51492 45726
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50428 45276 50484 45332
rect 50652 45218 50708 45220
rect 50652 45166 50654 45218
rect 50654 45166 50706 45218
rect 50706 45166 50708 45218
rect 50652 45164 50708 45166
rect 50428 44492 50484 44548
rect 51660 45500 51716 45556
rect 51548 45052 51604 45108
rect 48188 43596 48244 43652
rect 46396 42924 46452 42980
rect 47404 42978 47460 42980
rect 47404 42926 47406 42978
rect 47406 42926 47458 42978
rect 47458 42926 47460 42978
rect 47404 42924 47460 42926
rect 45836 41244 45892 41300
rect 46396 41804 46452 41860
rect 46508 41244 46564 41300
rect 47180 41244 47236 41300
rect 46844 40684 46900 40740
rect 46508 40572 46564 40628
rect 47180 40572 47236 40628
rect 49308 42476 49364 42532
rect 48748 41970 48804 41972
rect 48748 41918 48750 41970
rect 48750 41918 48802 41970
rect 48802 41918 48804 41970
rect 48748 41916 48804 41918
rect 49084 41916 49140 41972
rect 47964 40514 48020 40516
rect 47964 40462 47966 40514
rect 47966 40462 48018 40514
rect 48018 40462 48020 40514
rect 47964 40460 48020 40462
rect 78204 46396 78260 46452
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 50876 44828 50932 44884
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 51884 45948 51940 46004
rect 77644 45890 77700 45892
rect 77644 45838 77646 45890
rect 77646 45838 77698 45890
rect 77698 45838 77700 45890
rect 77644 45836 77700 45838
rect 77420 45778 77476 45780
rect 77420 45726 77422 45778
rect 77422 45726 77474 45778
rect 77474 45726 77476 45778
rect 77420 45724 77476 45726
rect 78204 45778 78260 45780
rect 78204 45726 78206 45778
rect 78206 45726 78258 45778
rect 78258 45726 78260 45778
rect 78204 45724 78260 45726
rect 52668 45612 52724 45668
rect 52108 45106 52164 45108
rect 52108 45054 52110 45106
rect 52110 45054 52162 45106
rect 52162 45054 52164 45106
rect 52108 45052 52164 45054
rect 52220 44156 52276 44212
rect 53340 44940 53396 44996
rect 54236 44994 54292 44996
rect 54236 44942 54238 44994
rect 54238 44942 54290 44994
rect 54290 44942 54292 44994
rect 54236 44940 54292 44942
rect 75404 44994 75460 44996
rect 75404 44942 75406 44994
rect 75406 44942 75458 44994
rect 75458 44942 75460 44994
rect 75404 44940 75460 44942
rect 77980 45052 78036 45108
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 50988 43708 51044 43764
rect 51212 43708 51268 43764
rect 51884 43708 51940 43764
rect 51884 42978 51940 42980
rect 51884 42926 51886 42978
rect 51886 42926 51938 42978
rect 51938 42926 51940 42978
rect 51884 42924 51940 42926
rect 50204 42476 50260 42532
rect 52892 44156 52948 44212
rect 78204 43762 78260 43764
rect 78204 43710 78206 43762
rect 78206 43710 78258 43762
rect 78258 43710 78260 43762
rect 78204 43708 78260 43710
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 52780 42978 52836 42980
rect 52780 42926 52782 42978
rect 52782 42926 52834 42978
rect 52834 42926 52836 42978
rect 52780 42924 52836 42926
rect 50428 42530 50484 42532
rect 50428 42478 50430 42530
rect 50430 42478 50482 42530
rect 50482 42478 50484 42530
rect 50428 42476 50484 42478
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50316 41916 50372 41972
rect 50652 41970 50708 41972
rect 50652 41918 50654 41970
rect 50654 41918 50706 41970
rect 50706 41918 50708 41970
rect 50652 41916 50708 41918
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 49532 40514 49588 40516
rect 49532 40462 49534 40514
rect 49534 40462 49586 40514
rect 49586 40462 49588 40514
rect 49532 40460 49588 40462
rect 51660 42476 51716 42532
rect 77980 42364 78036 42420
rect 53564 41858 53620 41860
rect 53564 41806 53566 41858
rect 53566 41806 53618 41858
rect 53618 41806 53620 41858
rect 53564 41804 53620 41806
rect 75292 41858 75348 41860
rect 75292 41806 75294 41858
rect 75294 41806 75346 41858
rect 75346 41806 75348 41858
rect 75292 41804 75348 41806
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 77868 41132 77924 41188
rect 77644 41074 77700 41076
rect 77644 41022 77646 41074
rect 77646 41022 77698 41074
rect 77698 41022 77700 41074
rect 77644 41020 77700 41022
rect 78204 41074 78260 41076
rect 78204 41022 78206 41074
rect 78206 41022 78258 41074
rect 78258 41022 78260 41074
rect 78204 41020 78260 41022
rect 77308 40908 77364 40964
rect 75292 40626 75348 40628
rect 75292 40574 75294 40626
rect 75294 40574 75346 40626
rect 75346 40574 75348 40626
rect 75292 40572 75348 40574
rect 78204 40348 78260 40404
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 44604 39564 44660 39620
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 42028 38668 42084 38724
rect 42364 38780 42420 38836
rect 40348 38556 40404 38612
rect 39788 37996 39844 38052
rect 39676 36988 39732 37044
rect 39564 36652 39620 36708
rect 39676 36482 39732 36484
rect 39676 36430 39678 36482
rect 39678 36430 39730 36482
rect 39730 36430 39732 36482
rect 39676 36428 39732 36430
rect 39340 36370 39396 36372
rect 39340 36318 39342 36370
rect 39342 36318 39394 36370
rect 39394 36318 39396 36370
rect 39340 36316 39396 36318
rect 39900 35420 39956 35476
rect 39900 34188 39956 34244
rect 41020 36706 41076 36708
rect 41020 36654 41022 36706
rect 41022 36654 41074 36706
rect 41074 36654 41076 36706
rect 41020 36652 41076 36654
rect 40684 36482 40740 36484
rect 40684 36430 40686 36482
rect 40686 36430 40738 36482
rect 40738 36430 40740 36482
rect 40684 36428 40740 36430
rect 40348 36316 40404 36372
rect 41356 36482 41412 36484
rect 41356 36430 41358 36482
rect 41358 36430 41410 36482
rect 41410 36430 41412 36482
rect 41356 36428 41412 36430
rect 41132 36316 41188 36372
rect 41132 35420 41188 35476
rect 40572 34860 40628 34916
rect 40012 33516 40068 33572
rect 40124 33906 40180 33908
rect 40124 33854 40126 33906
rect 40126 33854 40178 33906
rect 40178 33854 40180 33906
rect 40124 33852 40180 33854
rect 40908 34860 40964 34916
rect 40908 33852 40964 33908
rect 41580 36482 41636 36484
rect 41580 36430 41582 36482
rect 41582 36430 41634 36482
rect 41634 36430 41636 36482
rect 41580 36428 41636 36430
rect 41244 33852 41300 33908
rect 41356 34188 41412 34244
rect 42252 36428 42308 36484
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 78204 37660 78260 37716
rect 50764 37604 50820 37606
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 42364 36204 42420 36260
rect 42252 35532 42308 35588
rect 42140 34188 42196 34244
rect 40572 33458 40628 33460
rect 40572 33406 40574 33458
rect 40574 33406 40626 33458
rect 40626 33406 40628 33458
rect 40572 33404 40628 33406
rect 39228 33346 39284 33348
rect 39228 33294 39230 33346
rect 39230 33294 39282 33346
rect 39282 33294 39284 33346
rect 39228 33292 39284 33294
rect 40012 32450 40068 32452
rect 40012 32398 40014 32450
rect 40014 32398 40066 32450
rect 40066 32398 40068 32450
rect 40012 32396 40068 32398
rect 42364 34130 42420 34132
rect 42364 34078 42366 34130
rect 42366 34078 42418 34130
rect 42418 34078 42420 34130
rect 42364 34076 42420 34078
rect 41580 33404 41636 33460
rect 41580 32508 41636 32564
rect 39676 32002 39732 32004
rect 39676 31950 39678 32002
rect 39678 31950 39730 32002
rect 39730 31950 39732 32002
rect 39676 31948 39732 31950
rect 40348 31948 40404 32004
rect 39004 31554 39060 31556
rect 39004 31502 39006 31554
rect 39006 31502 39058 31554
rect 39058 31502 39060 31554
rect 39004 31500 39060 31502
rect 39116 30940 39172 30996
rect 39004 30380 39060 30436
rect 38556 30322 38612 30324
rect 38556 30270 38558 30322
rect 38558 30270 38610 30322
rect 38610 30270 38612 30322
rect 38556 30268 38612 30270
rect 38556 29650 38612 29652
rect 38556 29598 38558 29650
rect 38558 29598 38610 29650
rect 38610 29598 38612 29650
rect 38556 29596 38612 29598
rect 37884 29260 37940 29316
rect 37996 29372 38052 29428
rect 37772 29202 37828 29204
rect 37772 29150 37774 29202
rect 37774 29150 37826 29202
rect 37826 29150 37828 29202
rect 37772 29148 37828 29150
rect 37548 28476 37604 28532
rect 36540 27244 36596 27300
rect 37100 27244 37156 27300
rect 38220 28924 38276 28980
rect 41020 31666 41076 31668
rect 41020 31614 41022 31666
rect 41022 31614 41074 31666
rect 41074 31614 41076 31666
rect 41020 31612 41076 31614
rect 41020 31052 41076 31108
rect 41804 32396 41860 32452
rect 42140 33852 42196 33908
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 45388 35586 45444 35588
rect 45388 35534 45390 35586
rect 45390 35534 45442 35586
rect 45442 35534 45444 35586
rect 45388 35532 45444 35534
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 42588 34860 42644 34916
rect 43260 34860 43316 34916
rect 42700 34242 42756 34244
rect 42700 34190 42702 34242
rect 42702 34190 42754 34242
rect 42754 34190 42756 34242
rect 42700 34188 42756 34190
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 43036 34130 43092 34132
rect 43036 34078 43038 34130
rect 43038 34078 43090 34130
rect 43090 34078 43092 34130
rect 43036 34076 43092 34078
rect 42476 33404 42532 33460
rect 42252 33068 42308 33124
rect 41580 30994 41636 30996
rect 41580 30942 41582 30994
rect 41582 30942 41634 30994
rect 41634 30942 41636 30994
rect 41580 30940 41636 30942
rect 42140 31500 42196 31556
rect 39564 30882 39620 30884
rect 39564 30830 39566 30882
rect 39566 30830 39618 30882
rect 39618 30830 39620 30882
rect 39564 30828 39620 30830
rect 40460 30828 40516 30884
rect 39452 30380 39508 30436
rect 39788 29932 39844 29988
rect 39564 29260 39620 29316
rect 39452 29202 39508 29204
rect 39452 29150 39454 29202
rect 39454 29150 39506 29202
rect 39506 29150 39508 29202
rect 39452 29148 39508 29150
rect 39116 28476 39172 28532
rect 39900 29484 39956 29540
rect 42028 30434 42084 30436
rect 42028 30382 42030 30434
rect 42030 30382 42082 30434
rect 42082 30382 42084 30434
rect 42028 30380 42084 30382
rect 41020 30268 41076 30324
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 44044 33234 44100 33236
rect 44044 33182 44046 33234
rect 44046 33182 44098 33234
rect 44098 33182 44100 33234
rect 44044 33180 44100 33182
rect 45052 33180 45108 33236
rect 43484 31890 43540 31892
rect 43484 31838 43486 31890
rect 43486 31838 43538 31890
rect 43538 31838 43540 31890
rect 43484 31836 43540 31838
rect 43932 33122 43988 33124
rect 43932 33070 43934 33122
rect 43934 33070 43986 33122
rect 43986 33070 43988 33122
rect 43932 33068 43988 33070
rect 44156 32562 44212 32564
rect 44156 32510 44158 32562
rect 44158 32510 44210 32562
rect 44210 32510 44212 32562
rect 44156 32508 44212 32510
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 45052 32002 45108 32004
rect 45052 31950 45054 32002
rect 45054 31950 45106 32002
rect 45106 31950 45108 32002
rect 45052 31948 45108 31950
rect 42140 30268 42196 30324
rect 40684 29986 40740 29988
rect 40684 29934 40686 29986
rect 40686 29934 40738 29986
rect 40738 29934 40740 29986
rect 40684 29932 40740 29934
rect 43708 31612 43764 31668
rect 44828 31612 44884 31668
rect 45388 31554 45444 31556
rect 45388 31502 45390 31554
rect 45390 31502 45442 31554
rect 45442 31502 45444 31554
rect 45388 31500 45444 31502
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 43260 30380 43316 30436
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 78204 29708 78260 29764
rect 41020 29484 41076 29540
rect 39788 28924 39844 28980
rect 40348 28924 40404 28980
rect 39676 28028 39732 28084
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 78204 28924 78260 28980
rect 41020 28700 41076 28756
rect 40908 28082 40964 28084
rect 40908 28030 40910 28082
rect 40910 28030 40962 28082
rect 40962 28030 40964 28082
rect 40908 28028 40964 28030
rect 41916 28754 41972 28756
rect 41916 28702 41918 28754
rect 41918 28702 41970 28754
rect 41970 28702 41972 28754
rect 41916 28700 41972 28702
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 78204 28252 78260 28308
rect 50764 28196 50820 28198
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 78204 26908 78260 26964
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 78204 20242 78260 20244
rect 78204 20190 78206 20242
rect 78206 20190 78258 20242
rect 78258 20190 78260 20242
rect 78204 20188 78260 20190
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 28252 4172 28308 4228
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 78204 18844 78260 18900
rect 50764 18788 50820 18790
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 78428 16828 78484 16884
rect 78204 16156 78260 16212
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 78204 15484 78260 15540
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 36428 4172 36484 4228
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 79200 64596 80000 64624
rect 78194 64540 78204 64596
rect 78260 64540 80000 64596
rect 79200 64512 80000 64540
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 79200 60564 80000 60592
rect 78194 60508 78204 60564
rect 78260 60508 80000 60564
rect 79200 60480 80000 60508
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 79200 59892 80000 59920
rect 78194 59836 78204 59892
rect 78260 59836 80000 59892
rect 79200 59808 80000 59836
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 79200 57876 80000 57904
rect 78194 57820 78204 57876
rect 78260 57820 80000 57876
rect 79200 57792 80000 57820
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 79200 49812 80000 49840
rect 78194 49756 78204 49812
rect 78260 49756 80000 49812
rect 79200 49728 80000 49756
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 47842 49084 47852 49140
rect 47908 49084 49532 49140
rect 49588 49084 49598 49140
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 47618 48412 47628 48468
rect 47684 48412 48748 48468
rect 48804 48412 48814 48468
rect 47730 48300 47740 48356
rect 47796 48300 49756 48356
rect 49812 48300 49822 48356
rect 49074 48188 49084 48244
rect 49140 48188 49980 48244
rect 50036 48188 50046 48244
rect 49522 48076 49532 48132
rect 49588 48076 50540 48132
rect 50596 48076 50606 48132
rect 46274 47964 46284 48020
rect 46340 47964 47852 48020
rect 47908 47964 47918 48020
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 79200 47796 80000 47824
rect 77970 47740 77980 47796
rect 78036 47740 80000 47796
rect 79200 47712 80000 47740
rect 50530 47628 50540 47684
rect 50596 47628 51100 47684
rect 51156 47628 77868 47684
rect 77924 47628 77934 47684
rect 48738 47516 48748 47572
rect 48804 47516 49420 47572
rect 49476 47516 49486 47572
rect 48178 47404 48188 47460
rect 48244 47404 49196 47460
rect 49252 47404 49262 47460
rect 46834 47292 46844 47348
rect 46900 47292 47740 47348
rect 47796 47292 47806 47348
rect 51762 47292 51772 47348
rect 51828 47292 52668 47348
rect 52724 47292 52734 47348
rect 52882 47292 52892 47348
rect 52948 47292 53340 47348
rect 53396 47292 53676 47348
rect 53732 47292 75404 47348
rect 75460 47292 75470 47348
rect 29138 47180 29148 47236
rect 29204 47180 30492 47236
rect 30548 47180 30558 47236
rect 46274 47180 46284 47236
rect 46340 47180 46620 47236
rect 46676 47180 46686 47236
rect 48290 47180 48300 47236
rect 48356 47180 48636 47236
rect 48692 47180 48702 47236
rect 79200 47124 80000 47152
rect 30370 47068 30380 47124
rect 30436 47068 34636 47124
rect 34692 47068 34702 47124
rect 45826 47068 45836 47124
rect 45892 47068 46564 47124
rect 46722 47068 46732 47124
rect 46788 47068 47516 47124
rect 47572 47068 47582 47124
rect 77634 47068 77644 47124
rect 77700 47068 78204 47124
rect 78260 47068 80000 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 46508 47012 46564 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 79200 47040 80000 47068
rect 46508 46956 47460 47012
rect 47618 46956 47628 47012
rect 47684 46956 50204 47012
rect 50260 46956 50270 47012
rect 47404 46676 47460 46956
rect 47740 46844 49420 46900
rect 49476 46844 51100 46900
rect 51156 46844 51436 46900
rect 51492 46844 51502 46900
rect 47740 46676 47796 46844
rect 48290 46732 48300 46788
rect 48356 46732 49084 46788
rect 49140 46732 49150 46788
rect 50306 46732 50316 46788
rect 50372 46732 51884 46788
rect 51940 46732 51950 46788
rect 38546 46620 38556 46676
rect 38612 46620 42028 46676
rect 42084 46620 42094 46676
rect 45490 46620 45500 46676
rect 45556 46620 46396 46676
rect 46452 46620 46462 46676
rect 47394 46620 47404 46676
rect 47460 46620 47470 46676
rect 47730 46620 47740 46676
rect 47796 46620 47806 46676
rect 48514 46620 48524 46676
rect 48580 46620 48748 46676
rect 48804 46620 48814 46676
rect 49970 46620 49980 46676
rect 50036 46620 50876 46676
rect 50932 46620 50942 46676
rect 31266 46508 31276 46564
rect 31332 46508 31948 46564
rect 32004 46508 33068 46564
rect 33124 46508 33134 46564
rect 43026 46508 43036 46564
rect 43092 46508 46508 46564
rect 46564 46508 46574 46564
rect 47618 46508 47628 46564
rect 47684 46508 48636 46564
rect 48692 46508 48702 46564
rect 79200 46452 80000 46480
rect 47506 46396 47516 46452
rect 47572 46396 48860 46452
rect 48916 46396 49868 46452
rect 49924 46396 49934 46452
rect 78194 46396 78204 46452
rect 78260 46396 80000 46452
rect 79200 46368 80000 46396
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 49410 46172 49420 46228
rect 49476 46172 50988 46228
rect 51044 46172 51054 46228
rect 47170 46060 47180 46116
rect 47236 46060 49756 46116
rect 49812 46060 49822 46116
rect 50866 45948 50876 46004
rect 50932 45948 51884 46004
rect 51940 45948 51950 46004
rect 28466 45836 28476 45892
rect 28532 45836 29260 45892
rect 29316 45836 29326 45892
rect 32386 45836 32396 45892
rect 32452 45836 33292 45892
rect 33348 45836 33358 45892
rect 35410 45836 35420 45892
rect 35476 45836 36988 45892
rect 37044 45836 37054 45892
rect 50642 45836 50652 45892
rect 50708 45836 77644 45892
rect 77700 45836 77710 45892
rect 79200 45780 80000 45808
rect 35634 45724 35644 45780
rect 35700 45724 36428 45780
rect 36484 45724 36494 45780
rect 48626 45724 48636 45780
rect 48692 45724 50316 45780
rect 50372 45724 51436 45780
rect 51492 45724 51502 45780
rect 77410 45724 77420 45780
rect 77476 45724 78204 45780
rect 78260 45724 80000 45780
rect 79200 45696 80000 45724
rect 32162 45612 32172 45668
rect 32228 45612 33180 45668
rect 33236 45612 34076 45668
rect 34132 45612 35084 45668
rect 35140 45612 35150 45668
rect 48066 45612 48076 45668
rect 48132 45612 49420 45668
rect 49476 45612 49486 45668
rect 50372 45612 52668 45668
rect 52724 45612 52734 45668
rect 50372 45556 50428 45612
rect 46946 45500 46956 45556
rect 47012 45500 49868 45556
rect 49924 45500 50428 45556
rect 51650 45500 51660 45556
rect 51716 45500 51726 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 29922 45276 29932 45332
rect 29988 45276 31612 45332
rect 31668 45276 31678 45332
rect 33618 45276 33628 45332
rect 33684 45276 34412 45332
rect 34468 45276 35308 45332
rect 35364 45276 35374 45332
rect 39554 45276 39564 45332
rect 39620 45276 40348 45332
rect 40404 45276 41132 45332
rect 41188 45276 41198 45332
rect 47954 45276 47964 45332
rect 48020 45276 48860 45332
rect 48916 45276 50428 45332
rect 50484 45276 50494 45332
rect 51660 45220 51716 45500
rect 34290 45164 34300 45220
rect 34356 45164 34636 45220
rect 34692 45164 35532 45220
rect 35588 45164 35868 45220
rect 35924 45164 36316 45220
rect 36372 45164 36382 45220
rect 45266 45164 45276 45220
rect 45332 45164 46060 45220
rect 46116 45164 46126 45220
rect 50372 45164 50652 45220
rect 50708 45164 51716 45220
rect 33954 45052 33964 45108
rect 34020 45052 34748 45108
rect 34804 45052 34814 45108
rect 34962 45052 34972 45108
rect 35028 45052 36428 45108
rect 36484 45052 36494 45108
rect 45826 45052 45836 45108
rect 45892 45052 47068 45108
rect 47124 45052 47134 45108
rect 50372 44996 50428 45164
rect 43362 44940 43372 44996
rect 43428 44940 45948 44996
rect 46004 44940 46014 44996
rect 47842 44940 47852 44996
rect 47908 44940 48636 44996
rect 48692 44940 50428 44996
rect 50876 44884 50932 45164
rect 79200 45108 80000 45136
rect 51538 45052 51548 45108
rect 51604 45052 52108 45108
rect 52164 45052 52174 45108
rect 77970 45052 77980 45108
rect 78036 45052 80000 45108
rect 79200 45024 80000 45052
rect 53330 44940 53340 44996
rect 53396 44940 54236 44996
rect 54292 44940 75404 44996
rect 75460 44940 75470 44996
rect 30818 44828 30828 44884
rect 30884 44828 31724 44884
rect 31780 44828 31790 44884
rect 33842 44828 33852 44884
rect 33908 44828 34748 44884
rect 34804 44828 34814 44884
rect 38658 44828 38668 44884
rect 38724 44828 39788 44884
rect 39844 44828 39854 44884
rect 50866 44828 50876 44884
rect 50932 44828 50942 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 38994 44604 39004 44660
rect 39060 44604 39564 44660
rect 39620 44604 39630 44660
rect 35522 44492 35532 44548
rect 35588 44492 37212 44548
rect 37268 44492 39228 44548
rect 39284 44492 39294 44548
rect 49858 44492 49868 44548
rect 49924 44492 50428 44548
rect 50484 44492 50494 44548
rect 37874 44268 37884 44324
rect 37940 44268 39564 44324
rect 39620 44268 39630 44324
rect 42130 44156 42140 44212
rect 42196 44156 45388 44212
rect 45444 44156 45454 44212
rect 52210 44156 52220 44212
rect 52276 44156 52892 44212
rect 52948 44156 52958 44212
rect 44930 44044 44940 44100
rect 44996 44044 45724 44100
rect 45780 44044 45790 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 38434 43820 38444 43876
rect 38500 43820 38510 43876
rect 38444 43764 38500 43820
rect 38444 43708 39284 43764
rect 49746 43708 49756 43764
rect 49812 43708 50988 43764
rect 51044 43708 51212 43764
rect 51268 43708 51884 43764
rect 51940 43708 51950 43764
rect 78194 43708 78204 43764
rect 78260 43708 79268 43764
rect 39228 43652 39284 43708
rect 49756 43652 49812 43708
rect 30930 43596 30940 43652
rect 30996 43596 34300 43652
rect 34356 43596 34860 43652
rect 34916 43596 34926 43652
rect 38434 43596 38444 43652
rect 38500 43596 39172 43652
rect 39228 43596 39452 43652
rect 39508 43596 39518 43652
rect 48178 43596 48188 43652
rect 48244 43596 49812 43652
rect 39116 43540 39172 43596
rect 36306 43484 36316 43540
rect 36372 43484 38668 43540
rect 38724 43484 38734 43540
rect 39116 43484 39900 43540
rect 39956 43484 39966 43540
rect 79212 43428 79268 43708
rect 78988 43372 79268 43428
rect 29922 43260 29932 43316
rect 29988 43260 30716 43316
rect 30772 43260 30782 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 78988 43092 79044 43372
rect 79200 43092 80000 43120
rect 39554 43036 39564 43092
rect 39620 43036 40348 43092
rect 40404 43036 40414 43092
rect 78988 43036 80000 43092
rect 79200 43008 80000 43036
rect 45490 42924 45500 42980
rect 45556 42924 46396 42980
rect 46452 42924 47404 42980
rect 47460 42924 47470 42980
rect 51874 42924 51884 42980
rect 51940 42924 52780 42980
rect 52836 42924 52846 42980
rect 37202 42812 37212 42868
rect 37268 42812 38220 42868
rect 38276 42812 38286 42868
rect 32050 42700 32060 42756
rect 32116 42700 32508 42756
rect 32564 42700 33404 42756
rect 33460 42700 33470 42756
rect 36418 42700 36428 42756
rect 36484 42700 37436 42756
rect 37492 42700 38108 42756
rect 38164 42700 38174 42756
rect 33842 42476 33852 42532
rect 33908 42476 38892 42532
rect 38948 42476 38958 42532
rect 49298 42476 49308 42532
rect 49364 42476 50204 42532
rect 50260 42476 50428 42532
rect 50484 42476 51660 42532
rect 51716 42476 51726 42532
rect 79200 42420 80000 42448
rect 77970 42364 77980 42420
rect 78036 42364 80000 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 79200 42336 80000 42364
rect 38546 42140 38556 42196
rect 38612 42140 38622 42196
rect 38556 42084 38612 42140
rect 34962 42028 34972 42084
rect 35028 42028 37660 42084
rect 37716 42028 39116 42084
rect 39172 42028 39182 42084
rect 30818 41916 30828 41972
rect 30884 41916 31724 41972
rect 31780 41916 32396 41972
rect 32452 41916 33740 41972
rect 33796 41916 33806 41972
rect 38322 41916 38332 41972
rect 38388 41916 40796 41972
rect 40852 41916 40862 41972
rect 41122 41916 41132 41972
rect 41188 41916 41198 41972
rect 44930 41916 44940 41972
rect 44996 41916 45612 41972
rect 45668 41916 48748 41972
rect 48804 41916 48814 41972
rect 49074 41916 49084 41972
rect 49140 41916 50316 41972
rect 50372 41916 50652 41972
rect 50708 41916 50718 41972
rect 41132 41860 41188 41916
rect 28018 41804 28028 41860
rect 28084 41804 29260 41860
rect 29316 41804 29708 41860
rect 29764 41804 32956 41860
rect 33012 41804 33516 41860
rect 33572 41804 33582 41860
rect 38434 41804 38444 41860
rect 38500 41804 41188 41860
rect 45266 41804 45276 41860
rect 45332 41804 46396 41860
rect 46452 41804 46462 41860
rect 53554 41804 53564 41860
rect 53620 41804 75292 41860
rect 75348 41804 75358 41860
rect 31490 41692 31500 41748
rect 31556 41692 32060 41748
rect 32116 41692 32126 41748
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 28690 41356 28700 41412
rect 28756 41356 30604 41412
rect 30660 41356 30670 41412
rect 31154 41356 31164 41412
rect 31220 41356 32172 41412
rect 32228 41356 32238 41412
rect 38658 41356 38668 41412
rect 38724 41356 39452 41412
rect 39508 41356 39518 41412
rect 39890 41244 39900 41300
rect 39956 41244 41244 41300
rect 41300 41244 41310 41300
rect 43026 41244 43036 41300
rect 43092 41244 44156 41300
rect 44212 41244 45836 41300
rect 45892 41244 46508 41300
rect 46564 41244 47180 41300
rect 47236 41244 47246 41300
rect 38770 41132 38780 41188
rect 38836 41132 39564 41188
rect 39620 41132 39630 41188
rect 41458 41132 41468 41188
rect 41524 41132 42252 41188
rect 42308 41132 42812 41188
rect 42868 41132 43484 41188
rect 43540 41132 77868 41188
rect 77924 41132 77934 41188
rect 79200 41076 80000 41104
rect 35746 41020 35756 41076
rect 35812 41020 37436 41076
rect 37492 41020 41692 41076
rect 41748 41020 41758 41076
rect 77634 41020 77644 41076
rect 77700 41020 78204 41076
rect 78260 41020 78270 41076
rect 78428 41020 80000 41076
rect 78428 40964 78484 41020
rect 79200 40992 80000 41020
rect 43362 40908 43372 40964
rect 43428 40908 43932 40964
rect 43988 40908 43998 40964
rect 77298 40908 77308 40964
rect 77364 40908 78484 40964
rect 42018 40796 42028 40852
rect 42084 40796 42700 40852
rect 42756 40796 42766 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 37762 40572 37772 40628
rect 37828 40572 39228 40628
rect 39284 40572 39294 40628
rect 34626 40460 34636 40516
rect 34692 40460 35756 40516
rect 35812 40460 35822 40516
rect 37090 40460 37100 40516
rect 37156 40460 41020 40516
rect 41076 40460 41086 40516
rect 42028 40404 42084 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 46834 40684 46844 40740
rect 46900 40684 50428 40740
rect 50372 40628 50428 40684
rect 46498 40572 46508 40628
rect 46564 40572 47180 40628
rect 47236 40572 47246 40628
rect 50372 40572 75292 40628
rect 75348 40572 75358 40628
rect 47954 40460 47964 40516
rect 48020 40460 49532 40516
rect 49588 40460 49598 40516
rect 79200 40404 80000 40432
rect 31154 40348 31164 40404
rect 31220 40348 32060 40404
rect 32116 40348 32126 40404
rect 37874 40348 37884 40404
rect 37940 40348 42084 40404
rect 78194 40348 78204 40404
rect 78260 40348 80000 40404
rect 79200 40320 80000 40348
rect 30370 40236 30380 40292
rect 30436 40236 30716 40292
rect 30772 40236 34300 40292
rect 34356 40236 34366 40292
rect 31490 40012 31500 40068
rect 31556 40012 32060 40068
rect 32116 40012 32956 40068
rect 33012 40012 33022 40068
rect 38994 40012 39004 40068
rect 39060 40012 41132 40068
rect 41188 40012 41198 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 32386 39788 32396 39844
rect 32452 39788 32956 39844
rect 33012 39788 33022 39844
rect 32508 39732 32564 39788
rect 32498 39676 32508 39732
rect 32564 39676 32574 39732
rect 42018 39564 42028 39620
rect 42084 39564 42924 39620
rect 42980 39564 42990 39620
rect 43250 39564 43260 39620
rect 43316 39564 44604 39620
rect 44660 39564 44670 39620
rect 31826 39452 31836 39508
rect 31892 39452 32620 39508
rect 32676 39452 33180 39508
rect 33236 39452 33246 39508
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 41122 38780 41132 38836
rect 41188 38780 42364 38836
rect 42420 38780 42430 38836
rect 35522 38668 35532 38724
rect 35588 38668 36988 38724
rect 37044 38668 37054 38724
rect 40348 38668 42028 38724
rect 42084 38668 42094 38724
rect 40348 38612 40404 38668
rect 40338 38556 40348 38612
rect 40404 38556 40414 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 39218 38108 39228 38164
rect 39284 38108 39564 38164
rect 39620 38108 39630 38164
rect 30146 37996 30156 38052
rect 30212 37996 35084 38052
rect 35140 37996 35756 38052
rect 35812 37996 35822 38052
rect 35970 37996 35980 38052
rect 36036 37996 38556 38052
rect 38612 37996 39788 38052
rect 39844 37996 39854 38052
rect 34290 37884 34300 37940
rect 34356 37884 35420 37940
rect 35476 37884 35486 37940
rect 79200 37716 80000 37744
rect 78194 37660 78204 37716
rect 78260 37660 80000 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 79200 37632 80000 37660
rect 29138 36988 29148 37044
rect 29204 36988 33628 37044
rect 33684 36988 34748 37044
rect 34804 36988 34814 37044
rect 37986 36988 37996 37044
rect 38052 36988 39676 37044
rect 39732 36988 39742 37044
rect 36418 36876 36428 36932
rect 36484 36876 37324 36932
rect 37380 36876 38220 36932
rect 38276 36876 38668 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 38612 36820 38668 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 38612 36764 39116 36820
rect 39172 36764 39182 36820
rect 35522 36652 35532 36708
rect 35588 36652 36988 36708
rect 37044 36652 37054 36708
rect 39554 36652 39564 36708
rect 39620 36652 41020 36708
rect 41076 36652 41086 36708
rect 37650 36540 37660 36596
rect 37716 36540 38892 36596
rect 38948 36540 38958 36596
rect 39666 36428 39676 36484
rect 39732 36428 40684 36484
rect 40740 36428 41356 36484
rect 41412 36428 41422 36484
rect 41570 36428 41580 36484
rect 41636 36428 42252 36484
rect 42308 36428 42318 36484
rect 37314 36316 37324 36372
rect 37380 36316 38668 36372
rect 39330 36316 39340 36372
rect 39396 36316 40348 36372
rect 40404 36316 41132 36372
rect 41188 36316 41198 36372
rect 38612 36260 38668 36316
rect 31490 36204 31500 36260
rect 31556 36204 32172 36260
rect 32228 36204 32238 36260
rect 38612 36204 42364 36260
rect 42420 36204 42430 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 42242 35532 42252 35588
rect 42308 35532 45388 35588
rect 45444 35532 45454 35588
rect 39890 35420 39900 35476
rect 39956 35420 41132 35476
rect 41188 35420 41198 35476
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 38658 34860 38668 34916
rect 38724 34860 40572 34916
rect 40628 34860 40638 34916
rect 40898 34860 40908 34916
rect 40964 34860 42588 34916
rect 42644 34860 43260 34916
rect 43316 34860 43326 34916
rect 29922 34748 29932 34804
rect 29988 34748 31388 34804
rect 31444 34748 31454 34804
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 35634 34300 35644 34356
rect 35700 34300 36204 34356
rect 36260 34300 37100 34356
rect 37156 34300 37166 34356
rect 37426 34188 37436 34244
rect 37492 34188 38892 34244
rect 38948 34188 39900 34244
rect 39956 34188 39966 34244
rect 41346 34188 41356 34244
rect 41412 34188 42140 34244
rect 42196 34188 42700 34244
rect 42756 34188 42766 34244
rect 42354 34076 42364 34132
rect 42420 34076 43036 34132
rect 43092 34076 43102 34132
rect 31714 33852 31724 33908
rect 31780 33852 33852 33908
rect 33908 33852 35084 33908
rect 35140 33852 35150 33908
rect 40114 33852 40124 33908
rect 40180 33852 40908 33908
rect 40964 33852 40974 33908
rect 41234 33852 41244 33908
rect 41300 33852 42140 33908
rect 42196 33852 42206 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 38612 33516 40012 33572
rect 40068 33516 40078 33572
rect 38612 33460 38668 33516
rect 31266 33404 31276 33460
rect 31332 33404 33404 33460
rect 33460 33404 33470 33460
rect 34738 33404 34748 33460
rect 34804 33404 38668 33460
rect 40562 33404 40572 33460
rect 40628 33404 41580 33460
rect 41636 33404 42476 33460
rect 42532 33404 42542 33460
rect 32162 33292 32172 33348
rect 32228 33292 32238 33348
rect 32386 33292 32396 33348
rect 32452 33292 34972 33348
rect 35028 33292 35038 33348
rect 38322 33292 38332 33348
rect 38388 33292 39228 33348
rect 39284 33292 39294 33348
rect 32172 33236 32228 33292
rect 30930 33180 30940 33236
rect 30996 33180 31612 33236
rect 31668 33180 32228 33236
rect 44034 33180 44044 33236
rect 44100 33180 45052 33236
rect 45108 33180 45118 33236
rect 35970 33068 35980 33124
rect 36036 33068 37548 33124
rect 37604 33068 37614 33124
rect 42242 33068 42252 33124
rect 42308 33068 43932 33124
rect 43988 33068 43998 33124
rect 31938 32956 31948 33012
rect 32004 32956 34076 33012
rect 34132 32956 34142 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 32162 32844 32172 32900
rect 32228 32844 33964 32900
rect 34020 32844 34030 32900
rect 41570 32508 41580 32564
rect 41636 32508 44156 32564
rect 44212 32508 44222 32564
rect 40002 32396 40012 32452
rect 40068 32396 41804 32452
rect 41860 32396 41870 32452
rect 32386 32284 32396 32340
rect 32452 32284 33516 32340
rect 33572 32284 33582 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 38546 31948 38556 32004
rect 38612 31948 39676 32004
rect 39732 31948 39742 32004
rect 40338 31948 40348 32004
rect 40404 31948 45052 32004
rect 45108 31948 45118 32004
rect 43484 31892 43540 31948
rect 28130 31836 28140 31892
rect 28196 31836 29148 31892
rect 29204 31836 29214 31892
rect 31490 31836 31500 31892
rect 31556 31836 32172 31892
rect 32228 31836 32238 31892
rect 43474 31836 43484 31892
rect 43540 31836 43550 31892
rect 35970 31612 35980 31668
rect 36036 31612 37100 31668
rect 37156 31612 37166 31668
rect 41010 31612 41020 31668
rect 41076 31612 43708 31668
rect 43764 31612 44828 31668
rect 44884 31612 44894 31668
rect 28802 31500 28812 31556
rect 28868 31500 30604 31556
rect 30660 31500 30670 31556
rect 36082 31500 36092 31556
rect 36148 31500 38444 31556
rect 38500 31500 39004 31556
rect 39060 31500 39070 31556
rect 42130 31500 42140 31556
rect 42196 31500 45388 31556
rect 45444 31500 45454 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 32274 31164 32284 31220
rect 32340 31164 34300 31220
rect 34356 31164 37212 31220
rect 37268 31164 37278 31220
rect 36306 31052 36316 31108
rect 36372 31052 41020 31108
rect 41076 31052 41086 31108
rect 36754 30940 36764 30996
rect 36820 30940 39116 30996
rect 39172 30940 41580 30996
rect 41636 30940 41646 30996
rect 32498 30828 32508 30884
rect 32564 30828 33628 30884
rect 33684 30828 33694 30884
rect 39554 30828 39564 30884
rect 39620 30828 40460 30884
rect 40516 30828 40526 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 36194 30380 36204 30436
rect 36260 30380 36988 30436
rect 37044 30380 37054 30436
rect 38994 30380 39004 30436
rect 39060 30380 39452 30436
rect 39508 30380 42028 30436
rect 42084 30380 43260 30436
rect 43316 30380 43326 30436
rect 30482 30268 30492 30324
rect 30548 30268 31388 30324
rect 31444 30268 37548 30324
rect 37604 30268 37614 30324
rect 38546 30268 38556 30324
rect 38612 30268 41020 30324
rect 41076 30268 42140 30324
rect 42196 30268 42206 30324
rect 39778 29932 39788 29988
rect 39844 29932 40684 29988
rect 40740 29932 40750 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 78194 29708 78204 29764
rect 78260 29708 78270 29764
rect 78204 29652 78260 29708
rect 79200 29652 80000 29680
rect 36194 29596 36204 29652
rect 36260 29596 37100 29652
rect 37156 29596 37166 29652
rect 37762 29596 37772 29652
rect 37828 29596 38556 29652
rect 38612 29596 38622 29652
rect 78204 29596 80000 29652
rect 79200 29568 80000 29596
rect 39890 29484 39900 29540
rect 39956 29484 41020 29540
rect 41076 29484 41086 29540
rect 33506 29372 33516 29428
rect 33572 29372 35196 29428
rect 35252 29372 35262 29428
rect 36642 29372 36652 29428
rect 36708 29372 37996 29428
rect 38052 29372 38062 29428
rect 36418 29260 36428 29316
rect 36484 29260 37884 29316
rect 37940 29260 39564 29316
rect 39620 29260 39630 29316
rect 30146 29148 30156 29204
rect 30212 29148 31276 29204
rect 31332 29148 31342 29204
rect 32162 29148 32172 29204
rect 32228 29148 33740 29204
rect 33796 29148 33806 29204
rect 35410 29148 35420 29204
rect 35476 29148 36540 29204
rect 36596 29148 36606 29204
rect 37762 29148 37772 29204
rect 37828 29148 39452 29204
rect 39508 29148 39518 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 79200 28980 80000 29008
rect 38210 28924 38220 28980
rect 38276 28924 39788 28980
rect 39844 28924 40348 28980
rect 40404 28924 40414 28980
rect 78194 28924 78204 28980
rect 78260 28924 80000 28980
rect 79200 28896 80000 28924
rect 33842 28812 33852 28868
rect 33908 28812 35980 28868
rect 36036 28812 36046 28868
rect 41010 28700 41020 28756
rect 41076 28700 41916 28756
rect 41972 28700 41982 28756
rect 29362 28588 29372 28644
rect 29428 28588 32620 28644
rect 32676 28588 33964 28644
rect 34020 28588 34030 28644
rect 37538 28476 37548 28532
rect 37604 28476 39116 28532
rect 39172 28476 39182 28532
rect 79200 28308 80000 28336
rect 78194 28252 78204 28308
rect 78260 28252 80000 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 79200 28224 80000 28252
rect 39666 28028 39676 28084
rect 39732 28028 40908 28084
rect 40964 28028 40974 28084
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 36530 27244 36540 27300
rect 36596 27244 37100 27300
rect 37156 27244 37166 27300
rect 79200 26964 80000 26992
rect 78194 26908 78204 26964
rect 78260 26908 80000 26964
rect 79200 26880 80000 26908
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 78194 20188 78204 20244
rect 78260 20188 79268 20244
rect 79212 19796 79268 20188
rect 78988 19740 79268 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 78988 19572 79044 19740
rect 79200 19572 80000 19600
rect 78988 19516 80000 19572
rect 79200 19488 80000 19516
rect 79200 18900 80000 18928
rect 78194 18844 78204 18900
rect 78260 18844 80000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 79200 18816 80000 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 79200 16884 80000 16912
rect 78418 16828 78428 16884
rect 78484 16828 80000 16884
rect 79200 16800 80000 16828
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 79200 16212 80000 16240
rect 78194 16156 78204 16212
rect 78260 16156 80000 16212
rect 79200 16128 80000 16156
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 79200 15540 80000 15568
rect 78194 15484 78204 15540
rect 78260 15484 80000 15540
rect 79200 15456 80000 15484
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 28242 4172 28252 4228
rect 28308 4172 36428 4228
rect 36484 4172 36494 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38304 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _155_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _156_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34048 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32816 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _158_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _159_
timestamp 1698431365
transform 1 0 38752 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _160_
timestamp 1698431365
transform -1 0 42000 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40320 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38752 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _163_
timestamp 1698431365
transform 1 0 32256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _165_
timestamp 1698431365
transform -1 0 39312 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _166_
timestamp 1698431365
transform 1 0 36848 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _167_
timestamp 1698431365
transform 1 0 35504 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35840 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39200 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42448 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _171_
timestamp 1698431365
transform 1 0 37184 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39536 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _173_
timestamp 1698431365
transform -1 0 37520 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _174_
timestamp 1698431365
transform -1 0 37520 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _175_
timestamp 1698431365
transform -1 0 35952 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _176_
timestamp 1698431365
transform -1 0 35616 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _178_
timestamp 1698431365
transform -1 0 36176 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39088 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _180_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _181_
timestamp 1698431365
transform 1 0 36960 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _182_
timestamp 1698431365
transform 1 0 38752 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _183_
timestamp 1698431365
transform -1 0 41440 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39984 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _185_
timestamp 1698431365
transform -1 0 40544 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _186_
timestamp 1698431365
transform 1 0 41888 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _187_
timestamp 1698431365
transform -1 0 43120 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _188_
timestamp 1698431365
transform -1 0 42560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _189_
timestamp 1698431365
transform 1 0 39648 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _190_
timestamp 1698431365
transform -1 0 43456 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _191_
timestamp 1698431365
transform -1 0 43904 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _192_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1698431365
transform -1 0 44240 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _194_
timestamp 1698431365
transform -1 0 42672 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _195_
timestamp 1698431365
transform -1 0 36512 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _196_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38976 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1698431365
transform -1 0 37968 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _198_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43008 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _199_
timestamp 1698431365
transform 1 0 37520 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1698431365
transform -1 0 38976 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _201_
timestamp 1698431365
transform -1 0 41216 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41104 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _203_
timestamp 1698431365
transform -1 0 38304 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _204_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40208 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _205_
timestamp 1698431365
transform -1 0 35616 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _206_
timestamp 1698431365
transform -1 0 37520 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _207_
timestamp 1698431365
transform -1 0 36848 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _208_
timestamp 1698431365
transform -1 0 35840 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _209_
timestamp 1698431365
transform 1 0 35952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _210_
timestamp 1698431365
transform -1 0 38864 0 1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _211_
timestamp 1698431365
transform -1 0 34496 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _212_
timestamp 1698431365
transform -1 0 36400 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _213_
timestamp 1698431365
transform -1 0 34160 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _214_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _215_
timestamp 1698431365
transform -1 0 31808 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _216_
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _217_
timestamp 1698431365
transform 1 0 31808 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _218_
timestamp 1698431365
transform -1 0 33824 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _219_
timestamp 1698431365
transform 1 0 33264 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _220_
timestamp 1698431365
transform -1 0 31472 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _221_
timestamp 1698431365
transform -1 0 30912 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _222_
timestamp 1698431365
transform 1 0 32032 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _223_
timestamp 1698431365
transform -1 0 32704 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _224_
timestamp 1698431365
transform 1 0 31136 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _225_
timestamp 1698431365
transform 1 0 31136 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _226_
timestamp 1698431365
transform -1 0 32032 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _227_
timestamp 1698431365
transform -1 0 30576 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _228_
timestamp 1698431365
transform -1 0 34832 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _229_
timestamp 1698431365
transform 1 0 31472 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _230_
timestamp 1698431365
transform -1 0 32816 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _231_
timestamp 1698431365
transform -1 0 31920 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _232_
timestamp 1698431365
transform -1 0 31024 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _233_
timestamp 1698431365
transform -1 0 31920 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _234_
timestamp 1698431365
transform 1 0 31920 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _235_
timestamp 1698431365
transform -1 0 31360 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _236_
timestamp 1698431365
transform 1 0 32256 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _237_
timestamp 1698431365
transform 1 0 33824 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _238_
timestamp 1698431365
transform 1 0 31472 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _239_
timestamp 1698431365
transform -1 0 31472 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _240_
timestamp 1698431365
transform -1 0 31472 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _241_
timestamp 1698431365
transform -1 0 30800 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _242_
timestamp 1698431365
transform 1 0 31584 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _243_
timestamp 1698431365
transform 1 0 32928 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _244_
timestamp 1698431365
transform -1 0 34832 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _245_
timestamp 1698431365
transform -1 0 32368 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _246_
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _247_
timestamp 1698431365
transform 1 0 34272 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _248_
timestamp 1698431365
transform 1 0 34384 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _249_
timestamp 1698431365
transform 1 0 35056 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _250_
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _251_
timestamp 1698431365
transform -1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _252_
timestamp 1698431365
transform 1 0 34608 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _253_
timestamp 1698431365
transform 1 0 39424 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _254_
timestamp 1698431365
transform 1 0 39088 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _255_
timestamp 1698431365
transform -1 0 39088 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _256_
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _257_
timestamp 1698431365
transform 1 0 37968 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _258_
timestamp 1698431365
transform -1 0 39424 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _259_
timestamp 1698431365
transform 1 0 39200 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _260_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38864 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _261_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37072 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _262_
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _263_
timestamp 1698431365
transform -1 0 50848 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _264_
timestamp 1698431365
transform -1 0 51632 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _265_
timestamp 1698431365
transform -1 0 52192 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _266_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 51520 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _267_
timestamp 1698431365
transform 1 0 49616 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _268_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49728 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _269_
timestamp 1698431365
transform 1 0 49728 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _270_
timestamp 1698431365
transform 1 0 49952 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _271_
timestamp 1698431365
transform -1 0 50400 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _272_
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _273_
timestamp 1698431365
transform -1 0 52080 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _274_
timestamp 1698431365
transform -1 0 50624 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _275_
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _276_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 51296 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _277_
timestamp 1698431365
transform -1 0 47600 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _278_
timestamp 1698431365
transform -1 0 46928 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _279_
timestamp 1698431365
transform -1 0 46144 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _280_
timestamp 1698431365
transform -1 0 52976 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _281_
timestamp 1698431365
transform 1 0 50624 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _282_
timestamp 1698431365
transform 1 0 51296 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _283_
timestamp 1698431365
transform -1 0 48384 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _284_
timestamp 1698431365
transform -1 0 46704 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _285_
timestamp 1698431365
transform 1 0 45696 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _286_
timestamp 1698431365
transform 1 0 45360 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _287_
timestamp 1698431365
transform -1 0 49280 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _288_
timestamp 1698431365
transform -1 0 47824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _289_
timestamp 1698431365
transform 1 0 47824 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _290_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47264 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _291_
timestamp 1698431365
transform -1 0 49616 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _292_
timestamp 1698431365
transform -1 0 49728 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _293_
timestamp 1698431365
transform -1 0 49616 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _294_
timestamp 1698431365
transform -1 0 48496 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _295_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 47040 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _296_
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _297_
timestamp 1698431365
transform 1 0 47376 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _298_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _299_
timestamp 1698431365
transform -1 0 47376 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _300_
timestamp 1698431365
transform 1 0 45136 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _301_
timestamp 1698431365
transform 1 0 42560 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _302_
timestamp 1698431365
transform 1 0 47040 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _303_
timestamp 1698431365
transform 1 0 47488 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _304_
timestamp 1698431365
transform 1 0 46032 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _305_
timestamp 1698431365
transform 1 0 45472 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _306_
timestamp 1698431365
transform 1 0 42448 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _307_
timestamp 1698431365
transform 1 0 43680 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _308_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34608 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _309_
timestamp 1698431365
transform 1 0 33376 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _310_
timestamp 1698431365
transform -1 0 42448 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _311_
timestamp 1698431365
transform 1 0 38416 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _312_
timestamp 1698431365
transform 1 0 42336 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _313_
timestamp 1698431365
transform -1 0 44464 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _314_
timestamp 1698431365
transform 1 0 41440 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _315_
timestamp 1698431365
transform 1 0 36512 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _316_
timestamp 1698431365
transform 1 0 37296 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _317_
timestamp 1698431365
transform 1 0 38864 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _318_
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _319_
timestamp 1698431365
transform 1 0 32480 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _320_
timestamp 1698431365
transform 1 0 29232 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _321_
timestamp 1698431365
transform -1 0 34608 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _322_
timestamp 1698431365
transform 1 0 27888 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _323_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _324_
timestamp 1698431365
transform 1 0 28784 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _325_
timestamp 1698431365
transform 1 0 29456 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _326_
timestamp 1698431365
transform 1 0 27776 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _327_
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _328_
timestamp 1698431365
transform 1 0 28224 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _329_
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _330_
timestamp 1698431365
transform 1 0 32816 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _331_
timestamp 1698431365
transform -1 0 38640 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _332_
timestamp 1698431365
transform 1 0 38080 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _333_
timestamp 1698431365
transform -1 0 42224 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _334_
timestamp 1698431365
transform -1 0 38080 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _335_
timestamp 1698431365
transform 1 0 50512 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _336_
timestamp 1698431365
transform 1 0 51184 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _337_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _338_
timestamp 1698431365
transform 1 0 50624 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _339_
timestamp 1698431365
transform 1 0 42448 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _340_
timestamp 1698431365
transform 1 0 42112 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _341_
timestamp 1698431365
transform 1 0 41216 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _342_
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _343_
timestamp 1698431365
transform 1 0 46256 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _344_
timestamp 1698431365
transform 1 0 45136 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _345_
timestamp 1698431365
transform 1 0 42448 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__A1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41552 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__A1
timestamp 1698431365
transform -1 0 53536 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__A1
timestamp 1698431365
transform 1 0 53312 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__A1
timestamp 1698431365
transform -1 0 46368 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__I
timestamp 1698431365
transform -1 0 53424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__283__A1
timestamp 1698431365
transform 1 0 48832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__I
timestamp 1698431365
transform 1 0 49952 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__A1
timestamp 1698431365
transform -1 0 49504 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__A2
timestamp 1698431365
transform 1 0 50624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__A1
timestamp 1698431365
transform 1 0 51072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__I
timestamp 1698431365
transform -1 0 50624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A2
timestamp 1698431365
transform 1 0 50512 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__I
timestamp 1698431365
transform 1 0 43456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout11_I
timestamp 1698431365
transform -1 0 46368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 77728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 77504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 77728 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output4_I
timestamp 1698431365
transform 1 0 75264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output5_I
timestamp 1698431365
transform 1 0 75264 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output6_I
timestamp 1698431365
transform -1 0 75488 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output7_I
timestamp 1698431365
transform 1 0 50176 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output8_I
timestamp 1698431365
transform -1 0 75488 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1698431365
transform -1 0 38528 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1698431365
transform 1 0 37968 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1698431365
transform -1 0 38752 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1698431365
transform 1 0 38416 0 1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_13 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 77952 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_14
timestamp 1698431365
transform -1 0 58352 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_15
timestamp 1698431365
transform 1 0 77952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_16
timestamp 1698431365
transform -1 0 48944 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_17
timestamp 1698431365
transform -1 0 63056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_18
timestamp 1698431365
transform 1 0 77952 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_19
timestamp 1698431365
transform -1 0 59696 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_20
timestamp 1698431365
transform -1 0 51520 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_21
timestamp 1698431365
transform 1 0 77952 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_22
timestamp 1698431365
transform -1 0 67760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_23
timestamp 1698431365
transform 1 0 77952 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_24
timestamp 1698431365
transform -1 0 38864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_25
timestamp 1698431365
transform 1 0 77952 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_26
timestamp 1698431365
transform -1 0 26096 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_27
timestamp 1698431365
transform -1 0 30800 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_28
timestamp 1698431365
transform -1 0 34832 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_29
timestamp 1698431365
transform -1 0 59136 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_30
timestamp 1698431365
transform 1 0 77952 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_31
timestamp 1698431365
transform 1 0 77952 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_32
timestamp 1698431365
transform 1 0 77952 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_33
timestamp 1698431365
transform 1 0 77952 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_34
timestamp 1698431365
transform 1 0 77952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_35
timestamp 1698431365
transform 1 0 77952 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_36
timestamp 1698431365
transform -1 0 63728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_37
timestamp 1698431365
transform -1 0 61040 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_38
timestamp 1698431365
transform 1 0 77952 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_39
timestamp 1698431365
transform -1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_40
timestamp 1698431365
transform -1 0 59696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_41
timestamp 1698431365
transform -1 0 50624 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_42
timestamp 1698431365
transform -1 0 60368 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  control_system_43
timestamp 1698431365
transform -1 0 50288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  control_system_44 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 77952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  control_system_45
timestamp 1698431365
transform 1 0 77952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  control_system_46
timestamp 1698431365
transform -1 0 57008 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  control_system_47
timestamp 1698431365
transform -1 0 36288 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  control_system_48
timestamp 1698431365
transform -1 0 35504 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  control_system_49
timestamp 1698431365
transform 1 0 77952 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  control_system_50
timestamp 1698431365
transform 1 0 77952 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout9
timestamp 1698431365
transform -1 0 45136 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout10
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout11
timestamp 1698431365
transform -1 0 46144 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout12
timestamp 1698431365
transform 1 0 46144 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_290 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_298 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_300 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34944 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_324 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698431365
transform 1 0 38080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_330
timestamp 1698431365
transform 1 0 38304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_335
timestamp 1698431365
transform 1 0 38864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698431365
transform 1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_420
timestamp 1698431365
transform 1 0 48384 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_425
timestamp 1698431365
transform 1 0 48944 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_437
timestamp 1698431365
transform 1 0 50288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_441
timestamp 1698431365
transform 1 0 50736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_512
timestamp 1698431365
transform 1 0 58688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_516
timestamp 1698431365
transform 1 0 59136 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_521
timestamp 1698431365
transform 1 0 59696 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_537
timestamp 1698431365
transform 1 0 61488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_541
timestamp 1698431365
transform 1 0 61936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_543
timestamp 1698431365
transform 1 0 62160 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_546
timestamp 1698431365
transform 1 0 62496 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_551
timestamp 1698431365
transform 1 0 63056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_557
timestamp 1698431365
transform 1 0 63728 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_573
timestamp 1698431365
transform 1 0 65520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_577
timestamp 1698431365
transform 1 0 65968 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_580
timestamp 1698431365
transform 1 0 66304 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_588
timestamp 1698431365
transform 1 0 67200 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_593
timestamp 1698431365
transform 1 0 67760 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_609
timestamp 1698431365
transform 1 0 69552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_611
timestamp 1698431365
transform 1 0 69776 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_614
timestamp 1698431365
transform 1 0 70112 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_648
timestamp 1698431365
transform 1 0 73920 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_682
timestamp 1698431365
transform 1 0 77728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_686
timestamp 1698431365
transform 1 0 78176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698431365
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_556
timestamp 1698431365
transform 1 0 63616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_562
timestamp 1698431365
transform 1 0 64288 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_626
timestamp 1698431365
transform 1 0 71456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_632
timestamp 1698431365
transform 1 0 72128 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_664
timestamp 1698431365
transform 1 0 75712 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_680
timestamp 1698431365
transform 1 0 77504 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_521
timestamp 1698431365
transform 1 0 59696 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_527
timestamp 1698431365
transform 1 0 60368 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_591
timestamp 1698431365
transform 1 0 67536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_597
timestamp 1698431365
transform 1 0 68208 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_661
timestamp 1698431365
transform 1 0 75376 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_667
timestamp 1698431365
transform 1 0 76048 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_683
timestamp 1698431365
transform 1 0 77840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_687
timestamp 1698431365
transform 1 0 78288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_556
timestamp 1698431365
transform 1 0 63616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_562
timestamp 1698431365
transform 1 0 64288 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_626
timestamp 1698431365
transform 1 0 71456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_632
timestamp 1698431365
transform 1 0 72128 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_664
timestamp 1698431365
transform 1 0 75712 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_680
timestamp 1698431365
transform 1 0 77504 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_521
timestamp 1698431365
transform 1 0 59696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_527
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_591
timestamp 1698431365
transform 1 0 67536 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_597
timestamp 1698431365
transform 1 0 68208 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_661
timestamp 1698431365
transform 1 0 75376 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_667
timestamp 1698431365
transform 1 0 76048 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_683
timestamp 1698431365
transform 1 0 77840 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_687
timestamp 1698431365
transform 1 0 78288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_556
timestamp 1698431365
transform 1 0 63616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_562
timestamp 1698431365
transform 1 0 64288 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_626
timestamp 1698431365
transform 1 0 71456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_632
timestamp 1698431365
transform 1 0 72128 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_664
timestamp 1698431365
transform 1 0 75712 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_680
timestamp 1698431365
transform 1 0 77504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1698431365
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_527
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_591
timestamp 1698431365
transform 1 0 67536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_597
timestamp 1698431365
transform 1 0 68208 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_661
timestamp 1698431365
transform 1 0 75376 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_667
timestamp 1698431365
transform 1 0 76048 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_683
timestamp 1698431365
transform 1 0 77840 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_687
timestamp 1698431365
transform 1 0 78288 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_556
timestamp 1698431365
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_562
timestamp 1698431365
transform 1 0 64288 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_626
timestamp 1698431365
transform 1 0 71456 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_632
timestamp 1698431365
transform 1 0 72128 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_664
timestamp 1698431365
transform 1 0 75712 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_680
timestamp 1698431365
transform 1 0 77504 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_521
timestamp 1698431365
transform 1 0 59696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_591
timestamp 1698431365
transform 1 0 67536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_597
timestamp 1698431365
transform 1 0 68208 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_661
timestamp 1698431365
transform 1 0 75376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_667
timestamp 1698431365
transform 1 0 76048 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_683
timestamp 1698431365
transform 1 0 77840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_687
timestamp 1698431365
transform 1 0 78288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_556
timestamp 1698431365
transform 1 0 63616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_562
timestamp 1698431365
transform 1 0 64288 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_626
timestamp 1698431365
transform 1 0 71456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_632
timestamp 1698431365
transform 1 0 72128 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_664
timestamp 1698431365
transform 1 0 75712 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_680
timestamp 1698431365
transform 1 0 77504 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1698431365
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_527
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_591
timestamp 1698431365
transform 1 0 67536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_597
timestamp 1698431365
transform 1 0 68208 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_661
timestamp 1698431365
transform 1 0 75376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_667
timestamp 1698431365
transform 1 0 76048 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_683
timestamp 1698431365
transform 1 0 77840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_687
timestamp 1698431365
transform 1 0 78288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1698431365
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_562
timestamp 1698431365
transform 1 0 64288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_626
timestamp 1698431365
transform 1 0 71456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_632
timestamp 1698431365
transform 1 0 72128 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_664
timestamp 1698431365
transform 1 0 75712 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_680
timestamp 1698431365
transform 1 0 77504 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698431365
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698431365
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_527
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_591
timestamp 1698431365
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_597
timestamp 1698431365
transform 1 0 68208 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_661
timestamp 1698431365
transform 1 0 75376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_667
timestamp 1698431365
transform 1 0 76048 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_683
timestamp 1698431365
transform 1 0 77840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_687
timestamp 1698431365
transform 1 0 78288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698431365
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1698431365
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1698431365
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1698431365
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_632
timestamp 1698431365
transform 1 0 72128 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_664
timestamp 1698431365
transform 1 0 75712 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_680
timestamp 1698431365
transform 1 0 77504 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_521
timestamp 1698431365
transform 1 0 59696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1698431365
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_597
timestamp 1698431365
transform 1 0 68208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_661
timestamp 1698431365
transform 1 0 75376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_667
timestamp 1698431365
transform 1 0 76048 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_683
timestamp 1698431365
transform 1 0 77840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_687
timestamp 1698431365
transform 1 0 78288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698431365
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1698431365
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1698431365
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_632
timestamp 1698431365
transform 1 0 72128 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_664
timestamp 1698431365
transform 1 0 75712 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_680
timestamp 1698431365
transform 1 0 77504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1698431365
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1698431365
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1698431365
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1698431365
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_667
timestamp 1698431365
transform 1 0 76048 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_683
timestamp 1698431365
transform 1 0 77840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698431365
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_562
timestamp 1698431365
transform 1 0 64288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_626
timestamp 1698431365
transform 1 0 71456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_632
timestamp 1698431365
transform 1 0 72128 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_664
timestamp 1698431365
transform 1 0 75712 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_680
timestamp 1698431365
transform 1 0 77504 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_521
timestamp 1698431365
transform 1 0 59696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_527
timestamp 1698431365
transform 1 0 60368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_591
timestamp 1698431365
transform 1 0 67536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_597
timestamp 1698431365
transform 1 0 68208 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_661
timestamp 1698431365
transform 1 0 75376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_667
timestamp 1698431365
transform 1 0 76048 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_683
timestamp 1698431365
transform 1 0 77840 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698431365
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698431365
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_562
timestamp 1698431365
transform 1 0 64288 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_626
timestamp 1698431365
transform 1 0 71456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_632
timestamp 1698431365
transform 1 0 72128 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_664
timestamp 1698431365
transform 1 0 75712 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_680
timestamp 1698431365
transform 1 0 77504 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698431365
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_521
timestamp 1698431365
transform 1 0 59696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_527
timestamp 1698431365
transform 1 0 60368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_591
timestamp 1698431365
transform 1 0 67536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_597
timestamp 1698431365
transform 1 0 68208 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_661
timestamp 1698431365
transform 1 0 75376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_667
timestamp 1698431365
transform 1 0 76048 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_683
timestamp 1698431365
transform 1 0 77840 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698431365
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_556
timestamp 1698431365
transform 1 0 63616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_562
timestamp 1698431365
transform 1 0 64288 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_626
timestamp 1698431365
transform 1 0 71456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_632
timestamp 1698431365
transform 1 0 72128 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_664
timestamp 1698431365
transform 1 0 75712 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_680
timestamp 1698431365
transform 1 0 77504 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_381
timestamp 1698431365
transform 1 0 44016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_521
timestamp 1698431365
transform 1 0 59696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_527
timestamp 1698431365
transform 1 0 60368 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_591
timestamp 1698431365
transform 1 0 67536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_597
timestamp 1698431365
transform 1 0 68208 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_661
timestamp 1698431365
transform 1 0 75376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_667
timestamp 1698431365
transform 1 0 76048 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_683
timestamp 1698431365
transform 1 0 77840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_687
timestamp 1698431365
transform 1 0 78288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_556
timestamp 1698431365
transform 1 0 63616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_562
timestamp 1698431365
transform 1 0 64288 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_626
timestamp 1698431365
transform 1 0 71456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_632
timestamp 1698431365
transform 1 0 72128 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_664
timestamp 1698431365
transform 1 0 75712 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_680
timestamp 1698431365
transform 1 0 77504 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_521
timestamp 1698431365
transform 1 0 59696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_527
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_591
timestamp 1698431365
transform 1 0 67536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_597
timestamp 1698431365
transform 1 0 68208 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_661
timestamp 1698431365
transform 1 0 75376 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_667
timestamp 1698431365
transform 1 0 76048 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_683
timestamp 1698431365
transform 1 0 77840 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_687
timestamp 1698431365
transform 1 0 78288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698431365
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_556
timestamp 1698431365
transform 1 0 63616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_562
timestamp 1698431365
transform 1 0 64288 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_626
timestamp 1698431365
transform 1 0 71456 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_632
timestamp 1698431365
transform 1 0 72128 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_664
timestamp 1698431365
transform 1 0 75712 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_680
timestamp 1698431365
transform 1 0 77504 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698431365
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_521
timestamp 1698431365
transform 1 0 59696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_527
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_591
timestamp 1698431365
transform 1 0 67536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_597
timestamp 1698431365
transform 1 0 68208 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_661
timestamp 1698431365
transform 1 0 75376 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_667
timestamp 1698431365
transform 1 0 76048 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_683
timestamp 1698431365
transform 1 0 77840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_687
timestamp 1698431365
transform 1 0 78288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698431365
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_556
timestamp 1698431365
transform 1 0 63616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_562
timestamp 1698431365
transform 1 0 64288 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_626
timestamp 1698431365
transform 1 0 71456 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_632
timestamp 1698431365
transform 1 0 72128 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_664
timestamp 1698431365
transform 1 0 75712 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_680
timestamp 1698431365
transform 1 0 77504 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698431365
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_521
timestamp 1698431365
transform 1 0 59696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_527
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_591
timestamp 1698431365
transform 1 0 67536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_597
timestamp 1698431365
transform 1 0 68208 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_661
timestamp 1698431365
transform 1 0 75376 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_667
timestamp 1698431365
transform 1 0 76048 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_683
timestamp 1698431365
transform 1 0 77840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_687
timestamp 1698431365
transform 1 0 78288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698431365
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_556
timestamp 1698431365
transform 1 0 63616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_562
timestamp 1698431365
transform 1 0 64288 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_626
timestamp 1698431365
transform 1 0 71456 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_632
timestamp 1698431365
transform 1 0 72128 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_664
timestamp 1698431365
transform 1 0 75712 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_680
timestamp 1698431365
transform 1 0 77504 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_323
timestamp 1698431365
transform 1 0 37520 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_355
timestamp 1698431365
transform 1 0 41104 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_371
timestamp 1698431365
transform 1 0 42896 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_379
timestamp 1698431365
transform 1 0 43792 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_383
timestamp 1698431365
transform 1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_521
timestamp 1698431365
transform 1 0 59696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_527
timestamp 1698431365
transform 1 0 60368 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_591
timestamp 1698431365
transform 1 0 67536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_597
timestamp 1698431365
transform 1 0 68208 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_661
timestamp 1698431365
transform 1 0 75376 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_667
timestamp 1698431365
transform 1 0 76048 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_683
timestamp 1698431365
transform 1 0 77840 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_244
timestamp 1698431365
transform 1 0 28672 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_260
timestamp 1698431365
transform 1 0 30464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_264
timestamp 1698431365
transform 1 0 30912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_266
timestamp 1698431365
transform 1 0 31136 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_319
timestamp 1698431365
transform 1 0 37072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_356
timestamp 1698431365
transform 1 0 41216 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_556
timestamp 1698431365
transform 1 0 63616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_562
timestamp 1698431365
transform 1 0 64288 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_626
timestamp 1698431365
transform 1 0 71456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_632
timestamp 1698431365
transform 1 0 72128 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_664
timestamp 1698431365
transform 1 0 75712 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_680
timestamp 1698431365
transform 1 0 77504 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_313
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_364
timestamp 1698431365
transform 1 0 42112 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_380
timestamp 1698431365
transform 1 0 43904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_521
timestamp 1698431365
transform 1 0 59696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_527
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_591
timestamp 1698431365
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_597
timestamp 1698431365
transform 1 0 68208 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_661
timestamp 1698431365
transform 1 0 75376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_667
timestamp 1698431365
transform 1 0 76048 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_683
timestamp 1698431365
transform 1 0 77840 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_244
timestamp 1698431365
transform 1 0 28672 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_260
timestamp 1698431365
transform 1 0 30464 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_264
timestamp 1698431365
transform 1 0 30912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_272
timestamp 1698431365
transform 1 0 31808 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_284
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_293
timestamp 1698431365
transform 1 0 34160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_297
timestamp 1698431365
transform 1 0 34608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_299
timestamp 1698431365
transform 1 0 34832 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_308
timestamp 1698431365
transform 1 0 35840 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_321
timestamp 1698431365
transform 1 0 37296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_323
timestamp 1698431365
transform 1 0 37520 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_336
timestamp 1698431365
transform 1 0 38976 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_347
timestamp 1698431365
transform 1 0 40208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_556
timestamp 1698431365
transform 1 0 63616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_562
timestamp 1698431365
transform 1 0 64288 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_626
timestamp 1698431365
transform 1 0 71456 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_632
timestamp 1698431365
transform 1 0 72128 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_664
timestamp 1698431365
transform 1 0 75712 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_680
timestamp 1698431365
transform 1 0 77504 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_279
timestamp 1698431365
transform 1 0 32592 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_295
timestamp 1698431365
transform 1 0 34384 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_303
timestamp 1698431365
transform 1 0 35280 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_307
timestamp 1698431365
transform 1 0 35728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_313
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_321
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_323
timestamp 1698431365
transform 1 0 37520 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_336
timestamp 1698431365
transform 1 0 38976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_338
timestamp 1698431365
transform 1 0 39200 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_355
timestamp 1698431365
transform 1 0 41104 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_359
timestamp 1698431365
transform 1 0 41552 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_369
timestamp 1698431365
transform 1 0 42672 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698431365
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_521
timestamp 1698431365
transform 1 0 59696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_527
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_591
timestamp 1698431365
transform 1 0 67536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_597
timestamp 1698431365
transform 1 0 68208 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_661
timestamp 1698431365
transform 1 0 75376 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_667
timestamp 1698431365
transform 1 0 76048 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_683
timestamp 1698431365
transform 1 0 77840 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_236
timestamp 1698431365
transform 1 0 27776 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_266
timestamp 1698431365
transform 1 0 31136 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_270
timestamp 1698431365
transform 1 0 31584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_296
timestamp 1698431365
transform 1 0 34496 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_304
timestamp 1698431365
transform 1 0 35392 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_343
timestamp 1698431365
transform 1 0 39760 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_347
timestamp 1698431365
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_356
timestamp 1698431365
transform 1 0 41216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_387
timestamp 1698431365
transform 1 0 44688 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698431365
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_556
timestamp 1698431365
transform 1 0 63616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_562
timestamp 1698431365
transform 1 0 64288 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_626
timestamp 1698431365
transform 1 0 71456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_632
timestamp 1698431365
transform 1 0 72128 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_664
timestamp 1698431365
transform 1 0 75712 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_680
timestamp 1698431365
transform 1 0 77504 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_255
timestamp 1698431365
transform 1 0 29904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_257
timestamp 1698431365
transform 1 0 30128 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_264
timestamp 1698431365
transform 1 0 30912 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_297
timestamp 1698431365
transform 1 0 34608 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_339
timestamp 1698431365
transform 1 0 39312 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_380
timestamp 1698431365
transform 1 0 43904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_395
timestamp 1698431365
transform 1 0 45584 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_427
timestamp 1698431365
transform 1 0 49168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_443
timestamp 1698431365
transform 1 0 50960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698431365
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_521
timestamp 1698431365
transform 1 0 59696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_527
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_591
timestamp 1698431365
transform 1 0 67536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_597
timestamp 1698431365
transform 1 0 68208 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_661
timestamp 1698431365
transform 1 0 75376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_667
timestamp 1698431365
transform 1 0 76048 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_683
timestamp 1698431365
transform 1 0 77840 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_687
timestamp 1698431365
transform 1 0 78288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_244
timestamp 1698431365
transform 1 0 28672 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_252
timestamp 1698431365
transform 1 0 29568 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_269
timestamp 1698431365
transform 1 0 31472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_271
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_332
timestamp 1698431365
transform 1 0 38528 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_340
timestamp 1698431365
transform 1 0 39424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_385
timestamp 1698431365
transform 1 0 44464 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_417
timestamp 1698431365
transform 1 0 48048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_556
timestamp 1698431365
transform 1 0 63616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_562
timestamp 1698431365
transform 1 0 64288 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_626
timestamp 1698431365
transform 1 0 71456 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_632
timestamp 1698431365
transform 1 0 72128 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_664
timestamp 1698431365
transform 1 0 75712 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_680
timestamp 1698431365
transform 1 0 77504 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_263
timestamp 1698431365
transform 1 0 30800 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_265
timestamp 1698431365
transform 1 0 31024 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_285
timestamp 1698431365
transform 1 0 33264 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_289
timestamp 1698431365
transform 1 0 33712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_383
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698431365
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_521
timestamp 1698431365
transform 1 0 59696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_527
timestamp 1698431365
transform 1 0 60368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_591
timestamp 1698431365
transform 1 0 67536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_597
timestamp 1698431365
transform 1 0 68208 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_661
timestamp 1698431365
transform 1 0 75376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_667
timestamp 1698431365
transform 1 0 76048 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_683
timestamp 1698431365
transform 1 0 77840 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_687
timestamp 1698431365
transform 1 0 78288 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_244
timestamp 1698431365
transform 1 0 28672 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_260
timestamp 1698431365
transform 1 0 30464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_264
timestamp 1698431365
transform 1 0 30912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_274
timestamp 1698431365
transform 1 0 32032 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_284
timestamp 1698431365
transform 1 0 33152 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_293
timestamp 1698431365
transform 1 0 34160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_297
timestamp 1698431365
transform 1 0 34608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_299
timestamp 1698431365
transform 1 0 34832 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_306
timestamp 1698431365
transform 1 0 35616 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_324
timestamp 1698431365
transform 1 0 37632 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_340
timestamp 1698431365
transform 1 0 39424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_358
timestamp 1698431365
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_376
timestamp 1698431365
transform 1 0 43456 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_408
timestamp 1698431365
transform 1 0 47040 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_556
timestamp 1698431365
transform 1 0 63616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_562
timestamp 1698431365
transform 1 0 64288 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_626
timestamp 1698431365
transform 1 0 71456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_632
timestamp 1698431365
transform 1 0 72128 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_664
timestamp 1698431365
transform 1 0 75712 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_680
timestamp 1698431365
transform 1 0 77504 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_280
timestamp 1698431365
transform 1 0 32704 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_325
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_329
timestamp 1698431365
transform 1 0 38192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_360
timestamp 1698431365
transform 1 0 41664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_375
timestamp 1698431365
transform 1 0 43344 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698431365
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_521
timestamp 1698431365
transform 1 0 59696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_527
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_591
timestamp 1698431365
transform 1 0 67536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_597
timestamp 1698431365
transform 1 0 68208 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_661
timestamp 1698431365
transform 1 0 75376 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_667
timestamp 1698431365
transform 1 0 76048 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_683
timestamp 1698431365
transform 1 0 77840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_687
timestamp 1698431365
transform 1 0 78288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_360
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_364
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_395
timestamp 1698431365
transform 1 0 45584 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_411
timestamp 1698431365
transform 1 0 47376 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_556
timestamp 1698431365
transform 1 0 63616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_562
timestamp 1698431365
transform 1 0 64288 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_626
timestamp 1698431365
transform 1 0 71456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_632
timestamp 1698431365
transform 1 0 72128 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_664
timestamp 1698431365
transform 1 0 75712 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_680
timestamp 1698431365
transform 1 0 77504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_263
timestamp 1698431365
transform 1 0 30800 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_271
timestamp 1698431365
transform 1 0 31696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_273
timestamp 1698431365
transform 1 0 31920 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_280
timestamp 1698431365
transform 1 0 32704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_284
timestamp 1698431365
transform 1 0 33152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_323
timestamp 1698431365
transform 1 0 37520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_363
timestamp 1698431365
transform 1 0 42000 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_373
timestamp 1698431365
transform 1 0 43120 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_381
timestamp 1698431365
transform 1 0 44016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698431365
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_521
timestamp 1698431365
transform 1 0 59696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_527
timestamp 1698431365
transform 1 0 60368 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_591
timestamp 1698431365
transform 1 0 67536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_597
timestamp 1698431365
transform 1 0 68208 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_661
timestamp 1698431365
transform 1 0 75376 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_667
timestamp 1698431365
transform 1 0 76048 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_683
timestamp 1698431365
transform 1 0 77840 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_687
timestamp 1698431365
transform 1 0 78288 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_244
timestamp 1698431365
transform 1 0 28672 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_274
timestamp 1698431365
transform 1 0 32032 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_290
timestamp 1698431365
transform 1 0 33824 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_294
timestamp 1698431365
transform 1 0 34272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_296
timestamp 1698431365
transform 1 0 34496 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_334
timestamp 1698431365
transform 1 0 38752 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_556
timestamp 1698431365
transform 1 0 63616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_562
timestamp 1698431365
transform 1 0 64288 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_626
timestamp 1698431365
transform 1 0 71456 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_632
timestamp 1698431365
transform 1 0 72128 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_664
timestamp 1698431365
transform 1 0 75712 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_680
timestamp 1698431365
transform 1 0 77504 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_274
timestamp 1698431365
transform 1 0 32032 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_290
timestamp 1698431365
transform 1 0 33824 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_298
timestamp 1698431365
transform 1 0 34720 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_302
timestamp 1698431365
transform 1 0 35168 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_367
timestamp 1698431365
transform 1 0 42448 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_383
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_521
timestamp 1698431365
transform 1 0 59696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_527
timestamp 1698431365
transform 1 0 60368 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_591
timestamp 1698431365
transform 1 0 67536 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_597
timestamp 1698431365
transform 1 0 68208 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_661
timestamp 1698431365
transform 1 0 75376 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_667
timestamp 1698431365
transform 1 0 76048 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_683
timestamp 1698431365
transform 1 0 77840 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_244
timestamp 1698431365
transform 1 0 28672 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_248
timestamp 1698431365
transform 1 0 29120 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_250
timestamp 1698431365
transform 1 0 29344 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_298
timestamp 1698431365
transform 1 0 34720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_306
timestamp 1698431365
transform 1 0 35616 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_314
timestamp 1698431365
transform 1 0 36512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_316
timestamp 1698431365
transform 1 0 36736 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_323
timestamp 1698431365
transform 1 0 37520 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_330
timestamp 1698431365
transform 1 0 38304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_334
timestamp 1698431365
transform 1 0 38752 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_336
timestamp 1698431365
transform 1 0 38976 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_358
timestamp 1698431365
transform 1 0 41440 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_390
timestamp 1698431365
transform 1 0 45024 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_406
timestamp 1698431365
transform 1 0 46816 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_414
timestamp 1698431365
transform 1 0 47712 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_556
timestamp 1698431365
transform 1 0 63616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_562
timestamp 1698431365
transform 1 0 64288 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_626
timestamp 1698431365
transform 1 0 71456 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_632
timestamp 1698431365
transform 1 0 72128 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_664
timestamp 1698431365
transform 1 0 75712 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_680
timestamp 1698431365
transform 1 0 77504 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_287
timestamp 1698431365
transform 1 0 33488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_309
timestamp 1698431365
transform 1 0 35952 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_313
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_337
timestamp 1698431365
transform 1 0 39088 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_380
timestamp 1698431365
transform 1 0 43904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698431365
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_521
timestamp 1698431365
transform 1 0 59696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_527
timestamp 1698431365
transform 1 0 60368 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_591
timestamp 1698431365
transform 1 0 67536 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_597
timestamp 1698431365
transform 1 0 68208 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_661
timestamp 1698431365
transform 1 0 75376 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_667
timestamp 1698431365
transform 1 0 76048 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_683
timestamp 1698431365
transform 1 0 77840 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_687
timestamp 1698431365
transform 1 0 78288 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_244
timestamp 1698431365
transform 1 0 28672 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_260
timestamp 1698431365
transform 1 0 30464 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_268
timestamp 1698431365
transform 1 0 31360 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_277
timestamp 1698431365
transform 1 0 32368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_292
timestamp 1698431365
transform 1 0 34048 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_328
timestamp 1698431365
transform 1 0 38080 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_332
timestamp 1698431365
transform 1 0 38528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_334
timestamp 1698431365
transform 1 0 38752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_341
timestamp 1698431365
transform 1 0 39536 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_349
timestamp 1698431365
transform 1 0 40432 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_356
timestamp 1698431365
transform 1 0 41216 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_396
timestamp 1698431365
transform 1 0 45696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_398
timestamp 1698431365
transform 1 0 45920 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_405
timestamp 1698431365
transform 1 0 46704 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_409
timestamp 1698431365
transform 1 0 47152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_411
timestamp 1698431365
transform 1 0 47376 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_418
timestamp 1698431365
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_451
timestamp 1698431365
transform 1 0 51856 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_483
timestamp 1698431365
transform 1 0 55440 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_487
timestamp 1698431365
transform 1 0 55888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_489
timestamp 1698431365
transform 1 0 56112 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_556
timestamp 1698431365
transform 1 0 63616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_562
timestamp 1698431365
transform 1 0 64288 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_626
timestamp 1698431365
transform 1 0 71456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_632
timestamp 1698431365
transform 1 0 72128 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_648
timestamp 1698431365
transform 1 0 73920 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_656
timestamp 1698431365
transform 1 0 74816 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_255
timestamp 1698431365
transform 1 0 29904 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_259
timestamp 1698431365
transform 1 0 30352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_268
timestamp 1698431365
transform 1 0 31360 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_287
timestamp 1698431365
transform 1 0 33488 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_303
timestamp 1698431365
transform 1 0 35280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_319
timestamp 1698431365
transform 1 0 37072 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_326
timestamp 1698431365
transform 1 0 37856 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_335
timestamp 1698431365
transform 1 0 38864 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_365
timestamp 1698431365
transform 1 0 42224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_367
timestamp 1698431365
transform 1 0 42448 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_374
timestamp 1698431365
transform 1 0 43232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_391
timestamp 1698431365
transform 1 0 45136 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_393
timestamp 1698431365
transform 1 0 45360 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_400
timestamp 1698431365
transform 1 0 46144 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_430
timestamp 1698431365
transform 1 0 49504 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_446
timestamp 1698431365
transform 1 0 51296 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_454
timestamp 1698431365
transform 1 0 52192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_521
timestamp 1698431365
transform 1 0 59696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_527
timestamp 1698431365
transform 1 0 60368 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_591
timestamp 1698431365
transform 1 0 67536 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_597
timestamp 1698431365
transform 1 0 68208 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_661
timestamp 1698431365
transform 1 0 75376 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_667
timestamp 1698431365
transform 1 0 76048 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_675
timestamp 1698431365
transform 1 0 76944 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_679
timestamp 1698431365
transform 1 0 77392 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_228
timestamp 1698431365
transform 1 0 26880 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_360
timestamp 1698431365
transform 1 0 41664 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_376
timestamp 1698431365
transform 1 0 43456 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_384
timestamp 1698431365
transform 1 0 44352 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_428
timestamp 1698431365
transform 1 0 49280 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_436
timestamp 1698431365
transform 1 0 50176 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_438
timestamp 1698431365
transform 1 0 50400 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_468
timestamp 1698431365
transform 1 0 53760 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_484
timestamp 1698431365
transform 1 0 55552 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_488
timestamp 1698431365
transform 1 0 56000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_556
timestamp 1698431365
transform 1 0 63616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_562
timestamp 1698431365
transform 1 0 64288 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_626
timestamp 1698431365
transform 1 0 71456 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_632
timestamp 1698431365
transform 1 0 72128 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_648
timestamp 1698431365
transform 1 0 73920 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_656
timestamp 1698431365
transform 1 0 74816 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_276
timestamp 1698431365
transform 1 0 32256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_280
timestamp 1698431365
transform 1 0 32704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_291
timestamp 1698431365
transform 1 0 33936 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_307
timestamp 1698431365
transform 1 0 35728 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_391
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_393
timestamp 1698431365
transform 1 0 45360 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_416
timestamp 1698431365
transform 1 0 47936 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_432
timestamp 1698431365
transform 1 0 49728 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_453
timestamp 1698431365
transform 1 0 52080 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_462
timestamp 1698431365
transform 1 0 53088 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_466
timestamp 1698431365
transform 1 0 53536 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_498
timestamp 1698431365
transform 1 0 57120 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_514
timestamp 1698431365
transform 1 0 58912 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_522
timestamp 1698431365
transform 1 0 59808 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_524
timestamp 1698431365
transform 1 0 60032 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_527
timestamp 1698431365
transform 1 0 60368 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_591
timestamp 1698431365
transform 1 0 67536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_597
timestamp 1698431365
transform 1 0 68208 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_661
timestamp 1698431365
transform 1 0 75376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_667
timestamp 1698431365
transform 1 0 76048 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_683
timestamp 1698431365
transform 1 0 77840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_687
timestamp 1698431365
transform 1 0 78288 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_244
timestamp 1698431365
transform 1 0 28672 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_260
timestamp 1698431365
transform 1 0 30464 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_275
timestamp 1698431365
transform 1 0 32144 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_296
timestamp 1698431365
transform 1 0 34496 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_312
timestamp 1698431365
transform 1 0 36288 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_320
timestamp 1698431365
transform 1 0 37184 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_335
timestamp 1698431365
transform 1 0 38864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_337
timestamp 1698431365
transform 1 0 39088 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_360
timestamp 1698431365
transform 1 0 41664 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_364
timestamp 1698431365
transform 1 0 42112 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_366
timestamp 1698431365
transform 1 0 42336 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_396
timestamp 1698431365
transform 1 0 45696 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_402
timestamp 1698431365
transform 1 0 46368 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_418
timestamp 1698431365
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_438
timestamp 1698431365
transform 1 0 50400 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_448
timestamp 1698431365
transform 1 0 51520 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_480
timestamp 1698431365
transform 1 0 55104 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_488
timestamp 1698431365
transform 1 0 56000 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_556
timestamp 1698431365
transform 1 0 63616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_562
timestamp 1698431365
transform 1 0 64288 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_626
timestamp 1698431365
transform 1 0 71456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_632
timestamp 1698431365
transform 1 0 72128 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_664
timestamp 1698431365
transform 1 0 75712 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_680
timestamp 1698431365
transform 1 0 77504 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_279
timestamp 1698431365
transform 1 0 32592 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_306
timestamp 1698431365
transform 1 0 35616 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_325
timestamp 1698431365
transform 1 0 37744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_329
timestamp 1698431365
transform 1 0 38192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_331
timestamp 1698431365
transform 1 0 38416 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_346
timestamp 1698431365
transform 1 0 40096 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_354
timestamp 1698431365
transform 1 0 40992 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_399
timestamp 1698431365
transform 1 0 46032 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_405
timestamp 1698431365
transform 1 0 46704 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_421
timestamp 1698431365
transform 1 0 48496 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_429
timestamp 1698431365
transform 1 0 49392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_440
timestamp 1698431365
transform 1 0 50624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_442
timestamp 1698431365
transform 1 0 50848 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698431365
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_462
timestamp 1698431365
transform 1 0 53088 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_466
timestamp 1698431365
transform 1 0 53536 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_498
timestamp 1698431365
transform 1 0 57120 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_514
timestamp 1698431365
transform 1 0 58912 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_522
timestamp 1698431365
transform 1 0 59808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_524
timestamp 1698431365
transform 1 0 60032 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_527
timestamp 1698431365
transform 1 0 60368 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_591
timestamp 1698431365
transform 1 0 67536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_597
timestamp 1698431365
transform 1 0 68208 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_661
timestamp 1698431365
transform 1 0 75376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_667
timestamp 1698431365
transform 1 0 76048 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_683
timestamp 1698431365
transform 1 0 77840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_687
timestamp 1698431365
transform 1 0 78288 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_244
timestamp 1698431365
transform 1 0 28672 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_252
timestamp 1698431365
transform 1 0 29568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_277
timestamp 1698431365
transform 1 0 32368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_279
timestamp 1698431365
transform 1 0 32592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_296
timestamp 1698431365
transform 1 0 34496 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_343
timestamp 1698431365
transform 1 0 39760 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_347
timestamp 1698431365
transform 1 0 40208 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_384
timestamp 1698431365
transform 1 0 44352 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_392
timestamp 1698431365
transform 1 0 45248 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_404
timestamp 1698431365
transform 1 0 46592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_406
timestamp 1698431365
transform 1 0 46816 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_426
timestamp 1698431365
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_430
timestamp 1698431365
transform 1 0 49504 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_474
timestamp 1698431365
transform 1 0 54432 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_556
timestamp 1698431365
transform 1 0 63616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_562
timestamp 1698431365
transform 1 0 64288 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_626
timestamp 1698431365
transform 1 0 71456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_632
timestamp 1698431365
transform 1 0 72128 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_648
timestamp 1698431365
transform 1 0 73920 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_656
timestamp 1698431365
transform 1 0 74816 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_276
timestamp 1698431365
transform 1 0 32256 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_280
timestamp 1698431365
transform 1 0 32704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_290
timestamp 1698431365
transform 1 0 33824 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_299
timestamp 1698431365
transform 1 0 34832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_309
timestamp 1698431365
transform 1 0 35952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_313
timestamp 1698431365
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_325
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_327
timestamp 1698431365
transform 1 0 37968 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_357
timestamp 1698431365
transform 1 0 41328 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_373
timestamp 1698431365
transform 1 0 43120 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_381
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_403
timestamp 1698431365
transform 1 0 46480 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_431
timestamp 1698431365
transform 1 0 49616 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_438
timestamp 1698431365
transform 1 0 50400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_442
timestamp 1698431365
transform 1 0 50848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_454
timestamp 1698431365
transform 1 0 52192 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_521
timestamp 1698431365
transform 1 0 59696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_527
timestamp 1698431365
transform 1 0 60368 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_591
timestamp 1698431365
transform 1 0 67536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_597
timestamp 1698431365
transform 1 0 68208 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_661
timestamp 1698431365
transform 1 0 75376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_667
timestamp 1698431365
transform 1 0 76048 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_675
timestamp 1698431365
transform 1 0 76944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_677
timestamp 1698431365
transform 1 0 77168 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698431365
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_206
timestamp 1698431365
transform 1 0 24416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_228
timestamp 1698431365
transform 1 0 26880 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_236
timestamp 1698431365
transform 1 0 27776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_269
timestamp 1698431365
transform 1 0 31472 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_278
timestamp 1698431365
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_300
timestamp 1698431365
transform 1 0 34944 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_333
timestamp 1698431365
transform 1 0 38640 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_349
timestamp 1698431365
transform 1 0 40432 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_360
timestamp 1698431365
transform 1 0 41664 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_393
timestamp 1698431365
transform 1 0 45360 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_397
timestamp 1698431365
transform 1 0 45808 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_408
timestamp 1698431365
transform 1 0 47040 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_410
timestamp 1698431365
transform 1 0 47264 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_446
timestamp 1698431365
transform 1 0 51296 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_478
timestamp 1698431365
transform 1 0 54880 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698431365
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_556
timestamp 1698431365
transform 1 0 63616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_562
timestamp 1698431365
transform 1 0 64288 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_626
timestamp 1698431365
transform 1 0 71456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_632
timestamp 1698431365
transform 1 0 72128 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_664
timestamp 1698431365
transform 1 0 75712 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_680
timestamp 1698431365
transform 1 0 77504 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_241
timestamp 1698431365
transform 1 0 28336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_255
timestamp 1698431365
transform 1 0 29904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_263
timestamp 1698431365
transform 1 0 30800 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_279
timestamp 1698431365
transform 1 0 32592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_310
timestamp 1698431365
transform 1 0 36064 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698431365
transform 1 0 36512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_381
timestamp 1698431365
transform 1 0 44016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_391
timestamp 1698431365
transform 1 0 45136 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_397
timestamp 1698431365
transform 1 0 45808 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_399
timestamp 1698431365
transform 1 0 46032 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_431
timestamp 1698431365
transform 1 0 49616 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_437
timestamp 1698431365
transform 1 0 50288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_441
timestamp 1698431365
transform 1 0 50736 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_445
timestamp 1698431365
transform 1 0 51184 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698431365
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_461
timestamp 1698431365
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_465
timestamp 1698431365
transform 1 0 53424 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_497
timestamp 1698431365
transform 1 0 57008 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_513
timestamp 1698431365
transform 1 0 58800 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_521
timestamp 1698431365
transform 1 0 59696 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_527
timestamp 1698431365
transform 1 0 60368 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_591
timestamp 1698431365
transform 1 0 67536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_597
timestamp 1698431365
transform 1 0 68208 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_661
timestamp 1698431365
transform 1 0 75376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_667
timestamp 1698431365
transform 1 0 76048 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_675
timestamp 1698431365
transform 1 0 76944 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_679
timestamp 1698431365
transform 1 0 77392 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_346
timestamp 1698431365
transform 1 0 40096 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_384
timestamp 1698431365
transform 1 0 44352 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_392
timestamp 1698431365
transform 1 0 45248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_394
timestamp 1698431365
transform 1 0 45472 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_400
timestamp 1698431365
transform 1 0 46144 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_408
timestamp 1698431365
transform 1 0 47040 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_432
timestamp 1698431365
transform 1 0 49728 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_436
timestamp 1698431365
transform 1 0 50176 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_469
timestamp 1698431365
transform 1 0 53872 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_485
timestamp 1698431365
transform 1 0 55664 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_489
timestamp 1698431365
transform 1 0 56112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_556
timestamp 1698431365
transform 1 0 63616 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_562
timestamp 1698431365
transform 1 0 64288 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_626
timestamp 1698431365
transform 1 0 71456 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_632
timestamp 1698431365
transform 1 0 72128 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_648
timestamp 1698431365
transform 1 0 73920 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_656
timestamp 1698431365
transform 1 0 74816 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_241
timestamp 1698431365
transform 1 0 28336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_311
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_381
timestamp 1698431365
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_418
timestamp 1698431365
transform 1 0 48160 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_450
timestamp 1698431365
transform 1 0 51744 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_454
timestamp 1698431365
transform 1 0 52192 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_521
timestamp 1698431365
transform 1 0 59696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_527
timestamp 1698431365
transform 1 0 60368 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_591
timestamp 1698431365
transform 1 0 67536 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_597
timestamp 1698431365
transform 1 0 68208 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_661
timestamp 1698431365
transform 1 0 75376 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_667
timestamp 1698431365
transform 1 0 76048 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_683
timestamp 1698431365
transform 1 0 77840 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_687
timestamp 1698431365
transform 1 0 78288 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_346
timestamp 1698431365
transform 1 0 40096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698431365
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_486
timestamp 1698431365
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_556
timestamp 1698431365
transform 1 0 63616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_562
timestamp 1698431365
transform 1 0 64288 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_626
timestamp 1698431365
transform 1 0 71456 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_632
timestamp 1698431365
transform 1 0 72128 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_664
timestamp 1698431365
transform 1 0 75712 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_680
timestamp 1698431365
transform 1 0 77504 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_241
timestamp 1698431365
transform 1 0 28336 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_311
timestamp 1698431365
transform 1 0 36176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_381
timestamp 1698431365
transform 1 0 44016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_451
timestamp 1698431365
transform 1 0 51856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_521
timestamp 1698431365
transform 1 0 59696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_527
timestamp 1698431365
transform 1 0 60368 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_591
timestamp 1698431365
transform 1 0 67536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_597
timestamp 1698431365
transform 1 0 68208 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_661
timestamp 1698431365
transform 1 0 75376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_667
timestamp 1698431365
transform 1 0 76048 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_683
timestamp 1698431365
transform 1 0 77840 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698431365
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_276
timestamp 1698431365
transform 1 0 32256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_346
timestamp 1698431365
transform 1 0 40096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_416
timestamp 1698431365
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_486
timestamp 1698431365
transform 1 0 55776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_556
timestamp 1698431365
transform 1 0 63616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_562
timestamp 1698431365
transform 1 0 64288 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_626
timestamp 1698431365
transform 1 0 71456 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_632
timestamp 1698431365
transform 1 0 72128 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_664
timestamp 1698431365
transform 1 0 75712 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_680
timestamp 1698431365
transform 1 0 77504 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698431365
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_241
timestamp 1698431365
transform 1 0 28336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_311
timestamp 1698431365
transform 1 0 36176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_381
timestamp 1698431365
transform 1 0 44016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698431365
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_521
timestamp 1698431365
transform 1 0 59696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_527
timestamp 1698431365
transform 1 0 60368 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_591
timestamp 1698431365
transform 1 0 67536 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_597
timestamp 1698431365
transform 1 0 68208 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_661
timestamp 1698431365
transform 1 0 75376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_667
timestamp 1698431365
transform 1 0 76048 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_683
timestamp 1698431365
transform 1 0 77840 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_687
timestamp 1698431365
transform 1 0 78288 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698431365
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_276
timestamp 1698431365
transform 1 0 32256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_346
timestamp 1698431365
transform 1 0 40096 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_416
timestamp 1698431365
transform 1 0 47936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698431365
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_556
timestamp 1698431365
transform 1 0 63616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_562
timestamp 1698431365
transform 1 0 64288 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_626
timestamp 1698431365
transform 1 0 71456 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_632
timestamp 1698431365
transform 1 0 72128 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_664
timestamp 1698431365
transform 1 0 75712 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_680
timestamp 1698431365
transform 1 0 77504 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698431365
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_381
timestamp 1698431365
transform 1 0 44016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698431365
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_521
timestamp 1698431365
transform 1 0 59696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_527
timestamp 1698431365
transform 1 0 60368 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_591
timestamp 1698431365
transform 1 0 67536 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_597
timestamp 1698431365
transform 1 0 68208 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_661
timestamp 1698431365
transform 1 0 75376 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_667
timestamp 1698431365
transform 1 0 76048 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_683
timestamp 1698431365
transform 1 0 77840 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_687
timestamp 1698431365
transform 1 0 78288 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698431365
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_346
timestamp 1698431365
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_416
timestamp 1698431365
transform 1 0 47936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_556
timestamp 1698431365
transform 1 0 63616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_562
timestamp 1698431365
transform 1 0 64288 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_626
timestamp 1698431365
transform 1 0 71456 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_632
timestamp 1698431365
transform 1 0 72128 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_664
timestamp 1698431365
transform 1 0 75712 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_680
timestamp 1698431365
transform 1 0 77504 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698431365
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_241
timestamp 1698431365
transform 1 0 28336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_311
timestamp 1698431365
transform 1 0 36176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_381
timestamp 1698431365
transform 1 0 44016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_521
timestamp 1698431365
transform 1 0 59696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_527
timestamp 1698431365
transform 1 0 60368 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_591
timestamp 1698431365
transform 1 0 67536 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_597
timestamp 1698431365
transform 1 0 68208 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_661
timestamp 1698431365
transform 1 0 75376 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_667
timestamp 1698431365
transform 1 0 76048 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_683
timestamp 1698431365
transform 1 0 77840 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_687
timestamp 1698431365
transform 1 0 78288 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_66
timestamp 1698431365
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_136
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_276
timestamp 1698431365
transform 1 0 32256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_346
timestamp 1698431365
transform 1 0 40096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_416
timestamp 1698431365
transform 1 0 47936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_422
timestamp 1698431365
transform 1 0 48608 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_486
timestamp 1698431365
transform 1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_492
timestamp 1698431365
transform 1 0 56448 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_556
timestamp 1698431365
transform 1 0 63616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_562
timestamp 1698431365
transform 1 0 64288 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_626
timestamp 1698431365
transform 1 0 71456 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_632
timestamp 1698431365
transform 1 0 72128 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_664
timestamp 1698431365
transform 1 0 75712 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_680
timestamp 1698431365
transform 1 0 77504 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_37
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_101
timestamp 1698431365
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_171
timestamp 1698431365
transform 1 0 20496 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_177
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_241
timestamp 1698431365
transform 1 0 28336 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_247
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_311
timestamp 1698431365
transform 1 0 36176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_317
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_381
timestamp 1698431365
transform 1 0 44016 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_451
timestamp 1698431365
transform 1 0 51856 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_457
timestamp 1698431365
transform 1 0 52528 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_521
timestamp 1698431365
transform 1 0 59696 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_527
timestamp 1698431365
transform 1 0 60368 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_591
timestamp 1698431365
transform 1 0 67536 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_597
timestamp 1698431365
transform 1 0 68208 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_661
timestamp 1698431365
transform 1 0 75376 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_667
timestamp 1698431365
transform 1 0 76048 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_683
timestamp 1698431365
transform 1 0 77840 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_687
timestamp 1698431365
transform 1 0 78288 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_2
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_66
timestamp 1698431365
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_136
timestamp 1698431365
transform 1 0 16576 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_206
timestamp 1698431365
transform 1 0 24416 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_276
timestamp 1698431365
transform 1 0 32256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_346
timestamp 1698431365
transform 1 0 40096 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_416
timestamp 1698431365
transform 1 0 47936 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_422
timestamp 1698431365
transform 1 0 48608 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_486
timestamp 1698431365
transform 1 0 55776 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_492
timestamp 1698431365
transform 1 0 56448 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_556
timestamp 1698431365
transform 1 0 63616 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_562
timestamp 1698431365
transform 1 0 64288 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_626
timestamp 1698431365
transform 1 0 71456 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_632
timestamp 1698431365
transform 1 0 72128 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_664
timestamp 1698431365
transform 1 0 75712 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_680
timestamp 1698431365
transform 1 0 77504 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_2
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_101
timestamp 1698431365
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_171
timestamp 1698431365
transform 1 0 20496 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_241
timestamp 1698431365
transform 1 0 28336 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_311
timestamp 1698431365
transform 1 0 36176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_381
timestamp 1698431365
transform 1 0 44016 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_387
timestamp 1698431365
transform 1 0 44688 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_451
timestamp 1698431365
transform 1 0 51856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_457
timestamp 1698431365
transform 1 0 52528 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_521
timestamp 1698431365
transform 1 0 59696 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_527
timestamp 1698431365
transform 1 0 60368 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_591
timestamp 1698431365
transform 1 0 67536 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_597
timestamp 1698431365
transform 1 0 68208 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_661
timestamp 1698431365
transform 1 0 75376 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_667
timestamp 1698431365
transform 1 0 76048 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_683
timestamp 1698431365
transform 1 0 77840 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_66
timestamp 1698431365
transform 1 0 8736 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_136
timestamp 1698431365
transform 1 0 16576 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_206
timestamp 1698431365
transform 1 0 24416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_276
timestamp 1698431365
transform 1 0 32256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_282
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_346
timestamp 1698431365
transform 1 0 40096 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_352
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_416
timestamp 1698431365
transform 1 0 47936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_422
timestamp 1698431365
transform 1 0 48608 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_486
timestamp 1698431365
transform 1 0 55776 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_492
timestamp 1698431365
transform 1 0 56448 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_556
timestamp 1698431365
transform 1 0 63616 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_562
timestamp 1698431365
transform 1 0 64288 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_626
timestamp 1698431365
transform 1 0 71456 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_632
timestamp 1698431365
transform 1 0 72128 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_664
timestamp 1698431365
transform 1 0 75712 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_680
timestamp 1698431365
transform 1 0 77504 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_2
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_101
timestamp 1698431365
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_171
timestamp 1698431365
transform 1 0 20496 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_241
timestamp 1698431365
transform 1 0 28336 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_311
timestamp 1698431365
transform 1 0 36176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_381
timestamp 1698431365
transform 1 0 44016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_387
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_451
timestamp 1698431365
transform 1 0 51856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_457
timestamp 1698431365
transform 1 0 52528 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_521
timestamp 1698431365
transform 1 0 59696 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_527
timestamp 1698431365
transform 1 0 60368 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_591
timestamp 1698431365
transform 1 0 67536 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_597
timestamp 1698431365
transform 1 0 68208 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_661
timestamp 1698431365
transform 1 0 75376 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_667
timestamp 1698431365
transform 1 0 76048 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_683
timestamp 1698431365
transform 1 0 77840 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_2
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_66
timestamp 1698431365
transform 1 0 8736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_136
timestamp 1698431365
transform 1 0 16576 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_206
timestamp 1698431365
transform 1 0 24416 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_276
timestamp 1698431365
transform 1 0 32256 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_282
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_346
timestamp 1698431365
transform 1 0 40096 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_352
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_416
timestamp 1698431365
transform 1 0 47936 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_422
timestamp 1698431365
transform 1 0 48608 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_486
timestamp 1698431365
transform 1 0 55776 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_492
timestamp 1698431365
transform 1 0 56448 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_556
timestamp 1698431365
transform 1 0 63616 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_562
timestamp 1698431365
transform 1 0 64288 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_626
timestamp 1698431365
transform 1 0 71456 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_632
timestamp 1698431365
transform 1 0 72128 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_664
timestamp 1698431365
transform 1 0 75712 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_680
timestamp 1698431365
transform 1 0 77504 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1698431365
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_101
timestamp 1698431365
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_171
timestamp 1698431365
transform 1 0 20496 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_241
timestamp 1698431365
transform 1 0 28336 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_311
timestamp 1698431365
transform 1 0 36176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_381
timestamp 1698431365
transform 1 0 44016 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_387
timestamp 1698431365
transform 1 0 44688 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_451
timestamp 1698431365
transform 1 0 51856 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_457
timestamp 1698431365
transform 1 0 52528 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_521
timestamp 1698431365
transform 1 0 59696 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_527
timestamp 1698431365
transform 1 0 60368 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_591
timestamp 1698431365
transform 1 0 67536 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_597
timestamp 1698431365
transform 1 0 68208 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_661
timestamp 1698431365
transform 1 0 75376 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_667
timestamp 1698431365
transform 1 0 76048 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_683
timestamp 1698431365
transform 1 0 77840 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_687
timestamp 1698431365
transform 1 0 78288 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_2
timestamp 1698431365
transform 1 0 1568 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_66
timestamp 1698431365
transform 1 0 8736 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_136
timestamp 1698431365
transform 1 0 16576 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_206
timestamp 1698431365
transform 1 0 24416 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_276
timestamp 1698431365
transform 1 0 32256 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_346
timestamp 1698431365
transform 1 0 40096 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_352
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_416
timestamp 1698431365
transform 1 0 47936 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_422
timestamp 1698431365
transform 1 0 48608 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_486
timestamp 1698431365
transform 1 0 55776 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_492
timestamp 1698431365
transform 1 0 56448 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_556
timestamp 1698431365
transform 1 0 63616 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_562
timestamp 1698431365
transform 1 0 64288 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_626
timestamp 1698431365
transform 1 0 71456 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_632
timestamp 1698431365
transform 1 0 72128 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_664
timestamp 1698431365
transform 1 0 75712 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_680
timestamp 1698431365
transform 1 0 77504 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_2
timestamp 1698431365
transform 1 0 1568 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_101
timestamp 1698431365
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_171
timestamp 1698431365
transform 1 0 20496 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_241
timestamp 1698431365
transform 1 0 28336 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_311
timestamp 1698431365
transform 1 0 36176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_381
timestamp 1698431365
transform 1 0 44016 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_387
timestamp 1698431365
transform 1 0 44688 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_451
timestamp 1698431365
transform 1 0 51856 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_457
timestamp 1698431365
transform 1 0 52528 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_521
timestamp 1698431365
transform 1 0 59696 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_527
timestamp 1698431365
transform 1 0 60368 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_591
timestamp 1698431365
transform 1 0 67536 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_597
timestamp 1698431365
transform 1 0 68208 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_661
timestamp 1698431365
transform 1 0 75376 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_667
timestamp 1698431365
transform 1 0 76048 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_683
timestamp 1698431365
transform 1 0 77840 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_687
timestamp 1698431365
transform 1 0 78288 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_66
timestamp 1698431365
transform 1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_136
timestamp 1698431365
transform 1 0 16576 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_142
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_206
timestamp 1698431365
transform 1 0 24416 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_276
timestamp 1698431365
transform 1 0 32256 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_282
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_346
timestamp 1698431365
transform 1 0 40096 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_352
timestamp 1698431365
transform 1 0 40768 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_416
timestamp 1698431365
transform 1 0 47936 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_422
timestamp 1698431365
transform 1 0 48608 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_486
timestamp 1698431365
transform 1 0 55776 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_492
timestamp 1698431365
transform 1 0 56448 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_556
timestamp 1698431365
transform 1 0 63616 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_562
timestamp 1698431365
transform 1 0 64288 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_626
timestamp 1698431365
transform 1 0 71456 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_632
timestamp 1698431365
transform 1 0 72128 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_664
timestamp 1698431365
transform 1 0 75712 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_680
timestamp 1698431365
transform 1 0 77504 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_2
timestamp 1698431365
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_37
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_101
timestamp 1698431365
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_107
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_171
timestamp 1698431365
transform 1 0 20496 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_177
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_241
timestamp 1698431365
transform 1 0 28336 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_247
timestamp 1698431365
transform 1 0 29008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_311
timestamp 1698431365
transform 1 0 36176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_317
timestamp 1698431365
transform 1 0 36848 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_381
timestamp 1698431365
transform 1 0 44016 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_387
timestamp 1698431365
transform 1 0 44688 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_451
timestamp 1698431365
transform 1 0 51856 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_457
timestamp 1698431365
transform 1 0 52528 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_521
timestamp 1698431365
transform 1 0 59696 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_527
timestamp 1698431365
transform 1 0 60368 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_591
timestamp 1698431365
transform 1 0 67536 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_597
timestamp 1698431365
transform 1 0 68208 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_661
timestamp 1698431365
transform 1 0 75376 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_667
timestamp 1698431365
transform 1 0 76048 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_683
timestamp 1698431365
transform 1 0 77840 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_2
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_66
timestamp 1698431365
transform 1 0 8736 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_136
timestamp 1698431365
transform 1 0 16576 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_142
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_206
timestamp 1698431365
transform 1 0 24416 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_276
timestamp 1698431365
transform 1 0 32256 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_282
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_346
timestamp 1698431365
transform 1 0 40096 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_352
timestamp 1698431365
transform 1 0 40768 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_416
timestamp 1698431365
transform 1 0 47936 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_422
timestamp 1698431365
transform 1 0 48608 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_486
timestamp 1698431365
transform 1 0 55776 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_492
timestamp 1698431365
transform 1 0 56448 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_556
timestamp 1698431365
transform 1 0 63616 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_562
timestamp 1698431365
transform 1 0 64288 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_626
timestamp 1698431365
transform 1 0 71456 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_632
timestamp 1698431365
transform 1 0 72128 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_664
timestamp 1698431365
transform 1 0 75712 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_680
timestamp 1698431365
transform 1 0 77504 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_2
timestamp 1698431365
transform 1 0 1568 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_101
timestamp 1698431365
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_171
timestamp 1698431365
transform 1 0 20496 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_177
timestamp 1698431365
transform 1 0 21168 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_241
timestamp 1698431365
transform 1 0 28336 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_247
timestamp 1698431365
transform 1 0 29008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_311
timestamp 1698431365
transform 1 0 36176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_317
timestamp 1698431365
transform 1 0 36848 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_381
timestamp 1698431365
transform 1 0 44016 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_387
timestamp 1698431365
transform 1 0 44688 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_451
timestamp 1698431365
transform 1 0 51856 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_457
timestamp 1698431365
transform 1 0 52528 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_521
timestamp 1698431365
transform 1 0 59696 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_527
timestamp 1698431365
transform 1 0 60368 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_591
timestamp 1698431365
transform 1 0 67536 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_597
timestamp 1698431365
transform 1 0 68208 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_661
timestamp 1698431365
transform 1 0 75376 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_667
timestamp 1698431365
transform 1 0 76048 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_683
timestamp 1698431365
transform 1 0 77840 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_687
timestamp 1698431365
transform 1 0 78288 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_66
timestamp 1698431365
transform 1 0 8736 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_72
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_136
timestamp 1698431365
transform 1 0 16576 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_142
timestamp 1698431365
transform 1 0 17248 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_206
timestamp 1698431365
transform 1 0 24416 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_212
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_276
timestamp 1698431365
transform 1 0 32256 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_282
timestamp 1698431365
transform 1 0 32928 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_346
timestamp 1698431365
transform 1 0 40096 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_352
timestamp 1698431365
transform 1 0 40768 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_416
timestamp 1698431365
transform 1 0 47936 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_422
timestamp 1698431365
transform 1 0 48608 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_486
timestamp 1698431365
transform 1 0 55776 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_492
timestamp 1698431365
transform 1 0 56448 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_556
timestamp 1698431365
transform 1 0 63616 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_562
timestamp 1698431365
transform 1 0 64288 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_626
timestamp 1698431365
transform 1 0 71456 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_632
timestamp 1698431365
transform 1 0 72128 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_664
timestamp 1698431365
transform 1 0 75712 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_680
timestamp 1698431365
transform 1 0 77504 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_2
timestamp 1698431365
transform 1 0 1568 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1698431365
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_101
timestamp 1698431365
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_171
timestamp 1698431365
transform 1 0 20496 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_177
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_241
timestamp 1698431365
transform 1 0 28336 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_247
timestamp 1698431365
transform 1 0 29008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_311
timestamp 1698431365
transform 1 0 36176 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_317
timestamp 1698431365
transform 1 0 36848 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_381
timestamp 1698431365
transform 1 0 44016 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_387
timestamp 1698431365
transform 1 0 44688 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_451
timestamp 1698431365
transform 1 0 51856 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_457
timestamp 1698431365
transform 1 0 52528 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_521
timestamp 1698431365
transform 1 0 59696 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_527
timestamp 1698431365
transform 1 0 60368 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_591
timestamp 1698431365
transform 1 0 67536 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_597
timestamp 1698431365
transform 1 0 68208 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_661
timestamp 1698431365
transform 1 0 75376 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_667
timestamp 1698431365
transform 1 0 76048 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_683
timestamp 1698431365
transform 1 0 77840 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_687
timestamp 1698431365
transform 1 0 78288 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_2
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_66
timestamp 1698431365
transform 1 0 8736 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_72
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_136
timestamp 1698431365
transform 1 0 16576 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_142
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_206
timestamp 1698431365
transform 1 0 24416 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_212
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_276
timestamp 1698431365
transform 1 0 32256 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_282
timestamp 1698431365
transform 1 0 32928 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_346
timestamp 1698431365
transform 1 0 40096 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_352
timestamp 1698431365
transform 1 0 40768 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_416
timestamp 1698431365
transform 1 0 47936 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_422
timestamp 1698431365
transform 1 0 48608 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_486
timestamp 1698431365
transform 1 0 55776 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_492
timestamp 1698431365
transform 1 0 56448 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_556
timestamp 1698431365
transform 1 0 63616 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_562
timestamp 1698431365
transform 1 0 64288 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_626
timestamp 1698431365
transform 1 0 71456 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_632
timestamp 1698431365
transform 1 0 72128 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_664
timestamp 1698431365
transform 1 0 75712 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_680
timestamp 1698431365
transform 1 0 77504 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1698431365
transform 1 0 5152 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_101
timestamp 1698431365
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_107
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_171
timestamp 1698431365
transform 1 0 20496 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_241
timestamp 1698431365
transform 1 0 28336 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_247
timestamp 1698431365
transform 1 0 29008 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_311
timestamp 1698431365
transform 1 0 36176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_317
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_381
timestamp 1698431365
transform 1 0 44016 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_387
timestamp 1698431365
transform 1 0 44688 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_451
timestamp 1698431365
transform 1 0 51856 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_457
timestamp 1698431365
transform 1 0 52528 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_521
timestamp 1698431365
transform 1 0 59696 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_527
timestamp 1698431365
transform 1 0 60368 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_591
timestamp 1698431365
transform 1 0 67536 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_597
timestamp 1698431365
transform 1 0 68208 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_661
timestamp 1698431365
transform 1 0 75376 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_667
timestamp 1698431365
transform 1 0 76048 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_683
timestamp 1698431365
transform 1 0 77840 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_687
timestamp 1698431365
transform 1 0 78288 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_2
timestamp 1698431365
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_66
timestamp 1698431365
transform 1 0 8736 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_72
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_136
timestamp 1698431365
transform 1 0 16576 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_142
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_206
timestamp 1698431365
transform 1 0 24416 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_212
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_276
timestamp 1698431365
transform 1 0 32256 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_282
timestamp 1698431365
transform 1 0 32928 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_346
timestamp 1698431365
transform 1 0 40096 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_352
timestamp 1698431365
transform 1 0 40768 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_416
timestamp 1698431365
transform 1 0 47936 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_422
timestamp 1698431365
transform 1 0 48608 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_486
timestamp 1698431365
transform 1 0 55776 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_492
timestamp 1698431365
transform 1 0 56448 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_556
timestamp 1698431365
transform 1 0 63616 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_562
timestamp 1698431365
transform 1 0 64288 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_626
timestamp 1698431365
transform 1 0 71456 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_632
timestamp 1698431365
transform 1 0 72128 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_664
timestamp 1698431365
transform 1 0 75712 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_680
timestamp 1698431365
transform 1 0 77504 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_2
timestamp 1698431365
transform 1 0 1568 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_37
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_101
timestamp 1698431365
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_171
timestamp 1698431365
transform 1 0 20496 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_241
timestamp 1698431365
transform 1 0 28336 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_247
timestamp 1698431365
transform 1 0 29008 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_311
timestamp 1698431365
transform 1 0 36176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_317
timestamp 1698431365
transform 1 0 36848 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_381
timestamp 1698431365
transform 1 0 44016 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_387
timestamp 1698431365
transform 1 0 44688 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_451
timestamp 1698431365
transform 1 0 51856 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_457
timestamp 1698431365
transform 1 0 52528 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_521
timestamp 1698431365
transform 1 0 59696 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_527
timestamp 1698431365
transform 1 0 60368 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_591
timestamp 1698431365
transform 1 0 67536 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_597
timestamp 1698431365
transform 1 0 68208 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_661
timestamp 1698431365
transform 1 0 75376 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_667
timestamp 1698431365
transform 1 0 76048 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_683
timestamp 1698431365
transform 1 0 77840 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_687
timestamp 1698431365
transform 1 0 78288 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_66
timestamp 1698431365
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1698431365
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_206
timestamp 1698431365
transform 1 0 24416 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_276
timestamp 1698431365
transform 1 0 32256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_282
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_346
timestamp 1698431365
transform 1 0 40096 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_352
timestamp 1698431365
transform 1 0 40768 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_416
timestamp 1698431365
transform 1 0 47936 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_422
timestamp 1698431365
transform 1 0 48608 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_486
timestamp 1698431365
transform 1 0 55776 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_492
timestamp 1698431365
transform 1 0 56448 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_556
timestamp 1698431365
transform 1 0 63616 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_562
timestamp 1698431365
transform 1 0 64288 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_626
timestamp 1698431365
transform 1 0 71456 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_632
timestamp 1698431365
transform 1 0 72128 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_664
timestamp 1698431365
transform 1 0 75712 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_87_680
timestamp 1698431365
transform 1 0 77504 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_2
timestamp 1698431365
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698431365
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_101
timestamp 1698431365
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_171
timestamp 1698431365
transform 1 0 20496 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_241
timestamp 1698431365
transform 1 0 28336 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_247
timestamp 1698431365
transform 1 0 29008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_311
timestamp 1698431365
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_381
timestamp 1698431365
transform 1 0 44016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_387
timestamp 1698431365
transform 1 0 44688 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_451
timestamp 1698431365
transform 1 0 51856 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_457
timestamp 1698431365
transform 1 0 52528 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_521
timestamp 1698431365
transform 1 0 59696 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_527
timestamp 1698431365
transform 1 0 60368 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_591
timestamp 1698431365
transform 1 0 67536 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_597
timestamp 1698431365
transform 1 0 68208 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_661
timestamp 1698431365
transform 1 0 75376 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_667
timestamp 1698431365
transform 1 0 76048 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_683
timestamp 1698431365
transform 1 0 77840 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_687
timestamp 1698431365
transform 1 0 78288 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_2
timestamp 1698431365
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_66
timestamp 1698431365
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_72
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_136
timestamp 1698431365
transform 1 0 16576 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_206
timestamp 1698431365
transform 1 0 24416 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_276
timestamp 1698431365
transform 1 0 32256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_282
timestamp 1698431365
transform 1 0 32928 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_346
timestamp 1698431365
transform 1 0 40096 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_352
timestamp 1698431365
transform 1 0 40768 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_416
timestamp 1698431365
transform 1 0 47936 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_422
timestamp 1698431365
transform 1 0 48608 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_486
timestamp 1698431365
transform 1 0 55776 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_492
timestamp 1698431365
transform 1 0 56448 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_556
timestamp 1698431365
transform 1 0 63616 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_562
timestamp 1698431365
transform 1 0 64288 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_626
timestamp 1698431365
transform 1 0 71456 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_632
timestamp 1698431365
transform 1 0 72128 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_664
timestamp 1698431365
transform 1 0 75712 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_680
timestamp 1698431365
transform 1 0 77504 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_2
timestamp 1698431365
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1698431365
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_101
timestamp 1698431365
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_171
timestamp 1698431365
transform 1 0 20496 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_241
timestamp 1698431365
transform 1 0 28336 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_247
timestamp 1698431365
transform 1 0 29008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_311
timestamp 1698431365
transform 1 0 36176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_381
timestamp 1698431365
transform 1 0 44016 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_387
timestamp 1698431365
transform 1 0 44688 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_451
timestamp 1698431365
transform 1 0 51856 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_457
timestamp 1698431365
transform 1 0 52528 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_521
timestamp 1698431365
transform 1 0 59696 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_527
timestamp 1698431365
transform 1 0 60368 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_591
timestamp 1698431365
transform 1 0 67536 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_597
timestamp 1698431365
transform 1 0 68208 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_661
timestamp 1698431365
transform 1 0 75376 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_667
timestamp 1698431365
transform 1 0 76048 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_683
timestamp 1698431365
transform 1 0 77840 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_687
timestamp 1698431365
transform 1 0 78288 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_2
timestamp 1698431365
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_66
timestamp 1698431365
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_136
timestamp 1698431365
transform 1 0 16576 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_142
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_206
timestamp 1698431365
transform 1 0 24416 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_212
timestamp 1698431365
transform 1 0 25088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698431365
transform 1 0 32256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_282
timestamp 1698431365
transform 1 0 32928 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_346
timestamp 1698431365
transform 1 0 40096 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_352
timestamp 1698431365
transform 1 0 40768 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_416
timestamp 1698431365
transform 1 0 47936 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_422
timestamp 1698431365
transform 1 0 48608 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_486
timestamp 1698431365
transform 1 0 55776 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_492
timestamp 1698431365
transform 1 0 56448 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_556
timestamp 1698431365
transform 1 0 63616 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_562
timestamp 1698431365
transform 1 0 64288 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_626
timestamp 1698431365
transform 1 0 71456 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_632
timestamp 1698431365
transform 1 0 72128 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_664
timestamp 1698431365
transform 1 0 75712 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_680
timestamp 1698431365
transform 1 0 77504 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_2
timestamp 1698431365
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1698431365
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_101
timestamp 1698431365
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_171
timestamp 1698431365
transform 1 0 20496 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_177
timestamp 1698431365
transform 1 0 21168 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_241
timestamp 1698431365
transform 1 0 28336 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_247
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_311
timestamp 1698431365
transform 1 0 36176 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_317
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_381
timestamp 1698431365
transform 1 0 44016 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_387
timestamp 1698431365
transform 1 0 44688 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_419
timestamp 1698431365
transform 1 0 48272 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_435
timestamp 1698431365
transform 1 0 50064 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_438
timestamp 1698431365
transform 1 0 50400 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_454
timestamp 1698431365
transform 1 0 52192 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_457
timestamp 1698431365
transform 1 0 52528 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_521
timestamp 1698431365
transform 1 0 59696 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_527
timestamp 1698431365
transform 1 0 60368 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_591
timestamp 1698431365
transform 1 0 67536 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_597
timestamp 1698431365
transform 1 0 68208 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_661
timestamp 1698431365
transform 1 0 75376 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_667
timestamp 1698431365
transform 1 0 76048 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_683
timestamp 1698431365
transform 1 0 77840 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_687
timestamp 1698431365
transform 1 0 78288 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_2
timestamp 1698431365
transform 1 0 1568 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_36
timestamp 1698431365
transform 1 0 5376 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_70
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_104
timestamp 1698431365
transform 1 0 12992 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_138
timestamp 1698431365
transform 1 0 16800 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_172
timestamp 1698431365
transform 1 0 20608 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_206
timestamp 1698431365
transform 1 0 24416 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_214
timestamp 1698431365
transform 1 0 25312 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_216
timestamp 1698431365
transform 1 0 25536 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_221
timestamp 1698431365
transform 1 0 26096 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_237
timestamp 1698431365
transform 1 0 27888 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_240
timestamp 1698431365
transform 1 0 28224 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_256
timestamp 1698431365
transform 1 0 30016 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_258
timestamp 1698431365
transform 1 0 30240 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_263
timestamp 1698431365
transform 1 0 30800 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_271
timestamp 1698431365
transform 1 0 31696 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_274
timestamp 1698431365
transform 1 0 32032 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_290
timestamp 1698431365
transform 1 0 33824 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_294
timestamp 1698431365
transform 1 0 34272 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_299
timestamp 1698431365
transform 1 0 34832 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_305
timestamp 1698431365
transform 1 0 35504 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_312
timestamp 1698431365
transform 1 0 36288 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_328
timestamp 1698431365
transform 1 0 38080 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_336
timestamp 1698431365
transform 1 0 38976 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_342
timestamp 1698431365
transform 1 0 39648 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_376
timestamp 1698431365
transform 1 0 43456 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_440
timestamp 1698431365
transform 1 0 50624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_448
timestamp 1698431365
transform 1 0 51520 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_464
timestamp 1698431365
transform 1 0 53312 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_472
timestamp 1698431365
transform 1 0 54208 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_478
timestamp 1698431365
transform 1 0 54880 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_486
timestamp 1698431365
transform 1 0 55776 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_490
timestamp 1698431365
transform 1 0 56224 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_492
timestamp 1698431365
transform 1 0 56448 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_497
timestamp 1698431365
transform 1 0 57008 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_509
timestamp 1698431365
transform 1 0 58352 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_516
timestamp 1698431365
transform 1 0 59136 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_521
timestamp 1698431365
transform 1 0 59696 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_527
timestamp 1698431365
transform 1 0 60368 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_533
timestamp 1698431365
transform 1 0 61040 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_541
timestamp 1698431365
transform 1 0 61936 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_543
timestamp 1698431365
transform 1 0 62160 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_546
timestamp 1698431365
transform 1 0 62496 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_580
timestamp 1698431365
transform 1 0 66304 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_614
timestamp 1698431365
transform 1 0 70112 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_648
timestamp 1698431365
transform 1 0 73920 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_682
timestamp 1698431365
transform 1 0 77728 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_686
timestamp 1698431365
transform 1 0 78176 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform -1 0 78400 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698431365
transform -1 0 78400 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 78400 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 75488 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698431365
transform 1 0 75488 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698431365
transform 1 0 75488 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698431365
transform -1 0 50176 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698431365
transform 1 0 75488 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_136
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_137
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_138
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_139
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_140
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_141
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_142
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_143
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_144
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_145
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_146
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_147
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_148
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_149
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_150
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_151
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_152
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_153
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_154
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_155
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_156
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_157
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_158
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_159
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_160
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_161
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_162
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_163
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_164
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_165
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_166
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_167
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_168
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_169
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_170
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_171
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_172
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_173
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_174
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_175
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_176
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_177
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_178
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_179
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_180
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_181
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_182
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_183
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_184
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_185
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_186
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_187
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_188 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_189
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_190
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_191
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_192
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_193
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_194
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_195
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_196
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_197
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_198
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_199
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_200
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_201
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_202
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_203
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_204
timestamp 1698431365
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_205
timestamp 1698431365
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_206
timestamp 1698431365
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_207
timestamp 1698431365
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_208
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_209
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_210
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_211
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_212
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_213
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_214
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_215
timestamp 1698431365
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_216
timestamp 1698431365
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_217
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_218
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_219
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_220
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_221
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_222
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_223
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_224
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_225
timestamp 1698431365
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_226
timestamp 1698431365
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_227
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_228
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_229
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_230
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_231
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_232
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_233
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_234
timestamp 1698431365
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_235
timestamp 1698431365
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_236
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_237
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_238
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_239
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_240
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_241
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_242
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_243
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_244
timestamp 1698431365
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_245
timestamp 1698431365
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_246
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_247
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_248
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_249
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_250
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_251
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_252
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_253
timestamp 1698431365
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_254
timestamp 1698431365
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_255
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_256
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_257
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_258
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_259
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_260
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_261
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_262
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_263
timestamp 1698431365
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_264
timestamp 1698431365
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_265
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_266
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_267
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_268
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_269
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_270
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_271
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_272
timestamp 1698431365
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_273
timestamp 1698431365
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_274
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_275
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_276
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_277
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_278
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_279
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_280
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_281
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_282
timestamp 1698431365
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_283
timestamp 1698431365
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_284
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_285
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_286
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_287
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_288
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_289
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_290
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_291
timestamp 1698431365
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_292
timestamp 1698431365
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_293
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_294
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_295
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_296
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_297
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_298
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_299
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_300
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_301
timestamp 1698431365
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_302
timestamp 1698431365
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_303
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_304
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_305
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_306
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_307
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_308
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_309
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_310
timestamp 1698431365
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_311
timestamp 1698431365
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_312
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_313
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_314
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_315
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_316
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_317
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_318
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_319
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_320
timestamp 1698431365
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_321
timestamp 1698431365
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_322
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_323
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_324
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_325
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_326
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_327
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_328
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_329
timestamp 1698431365
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_330
timestamp 1698431365
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_331
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_332
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_333
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_334
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_335
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_336
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_337
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_338
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_339
timestamp 1698431365
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_340
timestamp 1698431365
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_341
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_342
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_343
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_344
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_345
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_346
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_347
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_348
timestamp 1698431365
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_349
timestamp 1698431365
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_350
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_351
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_352
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_353
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_354
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_355
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_356
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_357
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_358
timestamp 1698431365
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_359
timestamp 1698431365
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_360
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_361
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_362
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_363
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_364
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_365
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_366
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_367
timestamp 1698431365
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_368
timestamp 1698431365
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_369
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_370
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_371
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_372
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_373
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_374
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_375
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_376
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_377
timestamp 1698431365
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_378
timestamp 1698431365
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_379
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_380
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_381
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_382
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_383
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_384
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_385
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_386
timestamp 1698431365
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_387
timestamp 1698431365
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_388
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_389
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_390
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_391
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_392
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_393
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_394
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_395
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_396
timestamp 1698431365
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_397
timestamp 1698431365
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_398
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_399
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_400
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_401
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_402
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_403
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_404
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_405
timestamp 1698431365
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_406
timestamp 1698431365
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_407
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_408
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_409
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_410
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_411
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_412
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_413
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_414
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_415
timestamp 1698431365
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_416
timestamp 1698431365
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_417
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_418
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_419
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_420
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_421
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_422
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_423
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_424
timestamp 1698431365
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_425
timestamp 1698431365
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_426
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_427
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_428
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_429
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_430
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_431
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_432
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_433
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_434
timestamp 1698431365
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_435
timestamp 1698431365
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_436
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_437
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_438
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_439
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_440
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_441
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_442
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_443
timestamp 1698431365
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_444
timestamp 1698431365
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_445
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_446
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_447
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_448
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_449
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_450
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_451
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_452
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_453
timestamp 1698431365
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_454
timestamp 1698431365
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_455
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_456
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_457
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_458
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_459
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_460
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_461
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_462
timestamp 1698431365
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_463
timestamp 1698431365
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_464
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_465
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_466
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_467
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_468
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_469
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_470
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_471
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_472
timestamp 1698431365
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_473
timestamp 1698431365
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_474
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_475
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_476
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_477
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_478
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_479
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_480
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_481
timestamp 1698431365
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_482
timestamp 1698431365
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_483
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_484
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_485
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_486
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_487
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_488
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_489
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_490
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_491
timestamp 1698431365
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_492
timestamp 1698431365
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_493
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_494
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_495
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_496
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_497
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_498
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_499
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_500
timestamp 1698431365
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_501
timestamp 1698431365
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_502
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_503
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_504
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_505
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_506
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_507
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_508
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_509
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_510
timestamp 1698431365
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_511
timestamp 1698431365
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_512
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_513
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_514
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_515
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_516
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_517
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_518
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_519
timestamp 1698431365
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_520
timestamp 1698431365
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_521
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_522
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_523
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_524
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_525
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_526
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_527
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_528
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_529
timestamp 1698431365
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_530
timestamp 1698431365
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_531
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_532
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_533
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_534
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_535
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_536
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_537
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_538
timestamp 1698431365
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_539
timestamp 1698431365
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_540
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_541
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_542
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_543
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_544
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_545
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_546
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_547
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_548
timestamp 1698431365
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_549
timestamp 1698431365
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_550
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_551
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_552
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_553
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_554
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_555
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_556
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_557
timestamp 1698431365
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_558
timestamp 1698431365
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_559
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_560
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_561
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_562
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_563
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_564
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_565
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_566
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_567
timestamp 1698431365
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_568
timestamp 1698431365
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_569
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_570
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_571
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_572
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_573
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_574
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_575
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_576
timestamp 1698431365
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_577
timestamp 1698431365
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_578
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_579
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_580
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_581
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_582
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_583
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_584
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_585
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_586
timestamp 1698431365
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_587
timestamp 1698431365
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_588
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_589
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_590
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_591
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_592
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_593
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_594
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_595
timestamp 1698431365
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_596
timestamp 1698431365
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_597
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_598
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_599
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_600
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_601
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_602
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_603
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_604
timestamp 1698431365
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_605
timestamp 1698431365
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_606
timestamp 1698431365
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_607
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_608
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_609
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_610
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_611
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_612
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_613
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_614
timestamp 1698431365
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_615
timestamp 1698431365
transform 1 0 71904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_616
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_617
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_618
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_619
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_620
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_621
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_622
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_623
timestamp 1698431365
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_624
timestamp 1698431365
transform 1 0 67984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_625
timestamp 1698431365
transform 1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_626
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_627
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_628
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_629
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_630
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_631
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_632
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_633
timestamp 1698431365
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_634
timestamp 1698431365
transform 1 0 71904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_635
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_636
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_637
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_638
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_639
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_640
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_641
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_642
timestamp 1698431365
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_643
timestamp 1698431365
transform 1 0 67984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_644
timestamp 1698431365
transform 1 0 75824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_645
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_646
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_647
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_648
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_649
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_650
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_651
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_652
timestamp 1698431365
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_653
timestamp 1698431365
transform 1 0 71904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_654
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_655
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_656
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_657
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_658
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_659
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_660
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_661
timestamp 1698431365
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_662
timestamp 1698431365
transform 1 0 67984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_663
timestamp 1698431365
transform 1 0 75824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_664
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_665
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_666
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_667
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_668
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_669
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_670
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_671
timestamp 1698431365
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_672
timestamp 1698431365
transform 1 0 71904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_673
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_674
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_675
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_676
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_677
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_678
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_679
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_680
timestamp 1698431365
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_681
timestamp 1698431365
transform 1 0 67984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_682
timestamp 1698431365
transform 1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_683
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_684
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_685
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_686
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_687
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_688
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_689
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_690
timestamp 1698431365
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_691
timestamp 1698431365
transform 1 0 71904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_692
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_693
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_694
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_695
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_696
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_697
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_698
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_699
timestamp 1698431365
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_700
timestamp 1698431365
transform 1 0 67984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_701
timestamp 1698431365
transform 1 0 75824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_702
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_703
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_704
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_705
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_706
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_707
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_708
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_709
timestamp 1698431365
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_710
timestamp 1698431365
transform 1 0 71904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_711
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_712
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_713
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_714
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_715
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_716
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_717
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_718
timestamp 1698431365
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_719
timestamp 1698431365
transform 1 0 67984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_720
timestamp 1698431365
transform 1 0 75824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_721
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_722
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_723
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_724
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_725
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_726
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_727
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_728
timestamp 1698431365
transform 1 0 64064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_729
timestamp 1698431365
transform 1 0 71904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_730
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_731
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_732
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_733
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_734
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_735
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_736
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_737
timestamp 1698431365
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_738
timestamp 1698431365
transform 1 0 67984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_739
timestamp 1698431365
transform 1 0 75824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_740
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_741
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_742
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_743
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_744
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_745
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_746
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_747
timestamp 1698431365
transform 1 0 64064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_748
timestamp 1698431365
transform 1 0 71904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_749
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_750
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_751
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_752
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_753
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_754
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_755
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_756
timestamp 1698431365
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_757
timestamp 1698431365
transform 1 0 67984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_758
timestamp 1698431365
transform 1 0 75824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_759
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_760
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_761
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_762
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_763
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_764
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_765
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_766
timestamp 1698431365
transform 1 0 64064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_767
timestamp 1698431365
transform 1 0 71904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_768
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_769
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_770
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_771
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_772
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_773
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_774
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_775
timestamp 1698431365
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_776
timestamp 1698431365
transform 1 0 67984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_777
timestamp 1698431365
transform 1 0 75824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_778
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_779
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_780
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_781
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_782
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_783
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_784
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_785
timestamp 1698431365
transform 1 0 64064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_786
timestamp 1698431365
transform 1 0 71904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_787
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_788
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_789
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_790
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_791
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_792
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_793
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_794
timestamp 1698431365
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_795
timestamp 1698431365
transform 1 0 67984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_796
timestamp 1698431365
transform 1 0 75824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_797
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_798
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_799
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_800
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_801
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_802
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_803
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_804
timestamp 1698431365
transform 1 0 64064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_805
timestamp 1698431365
transform 1 0 71904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_806
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_807
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_808
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_809
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_810
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_811
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_812
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_813
timestamp 1698431365
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_814
timestamp 1698431365
transform 1 0 67984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_815
timestamp 1698431365
transform 1 0 75824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_816
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_817
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_818
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_819
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_820
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_821
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_822
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_823
timestamp 1698431365
transform 1 0 64064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_824
timestamp 1698431365
transform 1 0 71904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_825
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_826
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_827
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_828
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_829
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_830
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_831
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_832
timestamp 1698431365
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_833
timestamp 1698431365
transform 1 0 67984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_834
timestamp 1698431365
transform 1 0 75824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_835
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_836
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_837
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_838
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_839
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_840
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_841
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_842
timestamp 1698431365
transform 1 0 64064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_843
timestamp 1698431365
transform 1 0 71904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_844
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_845
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_846
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_847
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_848
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_849
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_850
timestamp 1698431365
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_851
timestamp 1698431365
transform 1 0 60144 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_852
timestamp 1698431365
transform 1 0 67984 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_853
timestamp 1698431365
transform 1 0 75824 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_854
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_855
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_856
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_857
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_858
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_859
timestamp 1698431365
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_860
timestamp 1698431365
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_861
timestamp 1698431365
transform 1 0 64064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_862
timestamp 1698431365
transform 1 0 71904 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_863
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_864
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_865
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_866
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_867
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_868
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_869
timestamp 1698431365
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_870
timestamp 1698431365
transform 1 0 60144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_871
timestamp 1698431365
transform 1 0 67984 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_872
timestamp 1698431365
transform 1 0 75824 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_873
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_874
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_875
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_876
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_877
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_878
timestamp 1698431365
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_879
timestamp 1698431365
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_880
timestamp 1698431365
transform 1 0 64064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_881
timestamp 1698431365
transform 1 0 71904 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_882
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_883
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_884
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_885
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_886
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_887
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_888
timestamp 1698431365
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_889
timestamp 1698431365
transform 1 0 60144 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_890
timestamp 1698431365
transform 1 0 67984 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_891
timestamp 1698431365
transform 1 0 75824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_892
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_893
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_894
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_895
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_896
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_897
timestamp 1698431365
transform 1 0 48384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_898
timestamp 1698431365
transform 1 0 56224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_899
timestamp 1698431365
transform 1 0 64064 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_900
timestamp 1698431365
transform 1 0 71904 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_901
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_902
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_903
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_904
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_905
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_906
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_907
timestamp 1698431365
transform 1 0 52304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_908
timestamp 1698431365
transform 1 0 60144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_909
timestamp 1698431365
transform 1 0 67984 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_910
timestamp 1698431365
transform 1 0 75824 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_911
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_912
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_913
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_914
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_915
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_916
timestamp 1698431365
transform 1 0 48384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_917
timestamp 1698431365
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_918
timestamp 1698431365
transform 1 0 64064 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_919
timestamp 1698431365
transform 1 0 71904 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_920
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_921
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_922
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_923
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_924
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_925
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_926
timestamp 1698431365
transform 1 0 52304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_927
timestamp 1698431365
transform 1 0 60144 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_928
timestamp 1698431365
transform 1 0 67984 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_929
timestamp 1698431365
transform 1 0 75824 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_930
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_931
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_932
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_933
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_934
timestamp 1698431365
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_935
timestamp 1698431365
transform 1 0 48384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_936
timestamp 1698431365
transform 1 0 56224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_937
timestamp 1698431365
transform 1 0 64064 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_938
timestamp 1698431365
transform 1 0 71904 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_939
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_940
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_941
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_942
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_943
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_944
timestamp 1698431365
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_945
timestamp 1698431365
transform 1 0 52304 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_946
timestamp 1698431365
transform 1 0 60144 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_947
timestamp 1698431365
transform 1 0 67984 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_948
timestamp 1698431365
transform 1 0 75824 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_949
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_950
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_951
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_952
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_953
timestamp 1698431365
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_954
timestamp 1698431365
transform 1 0 48384 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_955
timestamp 1698431365
transform 1 0 56224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_956
timestamp 1698431365
transform 1 0 64064 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_957
timestamp 1698431365
transform 1 0 71904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_958
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_959
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_960
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_961
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_962
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_963
timestamp 1698431365
transform 1 0 44464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_964
timestamp 1698431365
transform 1 0 52304 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_965
timestamp 1698431365
transform 1 0 60144 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_966
timestamp 1698431365
transform 1 0 67984 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_967
timestamp 1698431365
transform 1 0 75824 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_968
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_969
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_970
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_971
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_972
timestamp 1698431365
transform 1 0 40544 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_973
timestamp 1698431365
transform 1 0 48384 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_974
timestamp 1698431365
transform 1 0 56224 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_975
timestamp 1698431365
transform 1 0 64064 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_976
timestamp 1698431365
transform 1 0 71904 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_977
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_978
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_979
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_980
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_981
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_982
timestamp 1698431365
transform 1 0 44464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_983
timestamp 1698431365
transform 1 0 52304 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_984
timestamp 1698431365
transform 1 0 60144 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_985
timestamp 1698431365
transform 1 0 67984 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_986
timestamp 1698431365
transform 1 0 75824 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_987
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_988
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_989
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_990
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_991
timestamp 1698431365
transform 1 0 40544 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_992
timestamp 1698431365
transform 1 0 48384 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_993
timestamp 1698431365
transform 1 0 56224 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_994
timestamp 1698431365
transform 1 0 64064 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_995
timestamp 1698431365
transform 1 0 71904 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_996
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_997
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_998
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_999
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1000
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1001
timestamp 1698431365
transform 1 0 44464 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1002
timestamp 1698431365
transform 1 0 52304 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1003
timestamp 1698431365
transform 1 0 60144 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1004
timestamp 1698431365
transform 1 0 67984 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1005
timestamp 1698431365
transform 1 0 75824 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1006
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1007
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1008
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1009
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1010
timestamp 1698431365
transform 1 0 40544 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1011
timestamp 1698431365
transform 1 0 48384 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1012
timestamp 1698431365
transform 1 0 56224 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1013
timestamp 1698431365
transform 1 0 64064 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1014
timestamp 1698431365
transform 1 0 71904 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1015
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1016
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1017
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1018
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1019
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1020
timestamp 1698431365
transform 1 0 44464 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1021
timestamp 1698431365
transform 1 0 52304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1022
timestamp 1698431365
transform 1 0 60144 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1023
timestamp 1698431365
transform 1 0 67984 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1024
timestamp 1698431365
transform 1 0 75824 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1025
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1026
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1027
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1028
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1029
timestamp 1698431365
transform 1 0 40544 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1030
timestamp 1698431365
transform 1 0 48384 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1031
timestamp 1698431365
transform 1 0 56224 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1032
timestamp 1698431365
transform 1 0 64064 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1033
timestamp 1698431365
transform 1 0 71904 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1034
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1035
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1036
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1037
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1038
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1039
timestamp 1698431365
transform 1 0 44464 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1040
timestamp 1698431365
transform 1 0 52304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1041
timestamp 1698431365
transform 1 0 60144 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1042
timestamp 1698431365
transform 1 0 67984 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1043
timestamp 1698431365
transform 1 0 75824 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1044
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1045
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1046
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1047
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1048
timestamp 1698431365
transform 1 0 40544 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1049
timestamp 1698431365
transform 1 0 48384 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1050
timestamp 1698431365
transform 1 0 56224 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1051
timestamp 1698431365
transform 1 0 64064 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1052
timestamp 1698431365
transform 1 0 71904 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1053
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1054
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1055
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1056
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1057
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1058
timestamp 1698431365
transform 1 0 44464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1059
timestamp 1698431365
transform 1 0 52304 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1060
timestamp 1698431365
transform 1 0 60144 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1061
timestamp 1698431365
transform 1 0 67984 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1062
timestamp 1698431365
transform 1 0 75824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1063
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1064
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1065
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1066
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1067
timestamp 1698431365
transform 1 0 40544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1068
timestamp 1698431365
transform 1 0 48384 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1069
timestamp 1698431365
transform 1 0 56224 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1070
timestamp 1698431365
transform 1 0 64064 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1071
timestamp 1698431365
transform 1 0 71904 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1072
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1073
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1074
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1075
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1076
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1077
timestamp 1698431365
transform 1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1078
timestamp 1698431365
transform 1 0 52304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1079
timestamp 1698431365
transform 1 0 60144 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1080
timestamp 1698431365
transform 1 0 67984 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1081
timestamp 1698431365
transform 1 0 75824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1082
timestamp 1698431365
transform 1 0 5152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1083
timestamp 1698431365
transform 1 0 8960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1084
timestamp 1698431365
transform 1 0 12768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1085
timestamp 1698431365
transform 1 0 16576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1086
timestamp 1698431365
transform 1 0 20384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1087
timestamp 1698431365
transform 1 0 24192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1088
timestamp 1698431365
transform 1 0 28000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1089
timestamp 1698431365
transform 1 0 31808 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1090
timestamp 1698431365
transform 1 0 35616 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1091
timestamp 1698431365
transform 1 0 39424 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1092
timestamp 1698431365
transform 1 0 43232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1093
timestamp 1698431365
transform 1 0 47040 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1094
timestamp 1698431365
transform 1 0 50848 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1095
timestamp 1698431365
transform 1 0 54656 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1096
timestamp 1698431365
transform 1 0 58464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1097
timestamp 1698431365
transform 1 0 62272 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1098
timestamp 1698431365
transform 1 0 66080 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1099
timestamp 1698431365
transform 1 0 69888 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1100
timestamp 1698431365
transform 1 0 73696 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1101
timestamp 1698431365
transform 1 0 77504 0 -1 76832
box -86 -86 310 870
<< labels >>
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 79200 40992 80000 41104 0 FreeSans 448 0 0 0 clk_s
port 1 nsew signal tristate
flabel metal3 s 79200 47040 80000 47152 0 FreeSans 448 0 0 0 dir
port 2 nsew signal input
flabel metal3 s 79200 45696 80000 45808 0 FreeSans 448 0 0 0 enable
port 3 nsew signal input
flabel metal3 s 79200 26880 80000 26992 0 FreeSans 448 0 0 0 io_oeb[0]
port 4 nsew signal tristate
flabel metal2 s 48384 0 48496 800 0 FreeSans 448 90 0 0 io_oeb[10]
port 5 nsew signal tristate
flabel metal2 s 62496 0 62608 800 0 FreeSans 448 90 0 0 io_oeb[11]
port 6 nsew signal tristate
flabel metal3 s 79200 49728 80000 49840 0 FreeSans 448 0 0 0 io_oeb[12]
port 7 nsew signal tristate
flabel metal2 s 59136 79200 59248 80000 0 FreeSans 448 90 0 0 io_oeb[13]
port 8 nsew signal tristate
flabel metal2 s 50400 79200 50512 80000 0 FreeSans 448 90 0 0 io_oeb[14]
port 9 nsew signal tristate
flabel metal3 s 79200 28896 80000 29008 0 FreeSans 448 0 0 0 io_oeb[15]
port 10 nsew signal tristate
flabel metal2 s 67200 0 67312 800 0 FreeSans 448 90 0 0 io_oeb[16]
port 11 nsew signal tristate
flabel metal3 s 79200 16800 80000 16912 0 FreeSans 448 0 0 0 io_oeb[17]
port 12 nsew signal tristate
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 io_oeb[18]
port 13 nsew signal tristate
flabel metal3 s 79200 43008 80000 43120 0 FreeSans 448 0 0 0 io_oeb[19]
port 14 nsew signal tristate
flabel metal3 s 79200 29568 80000 29680 0 FreeSans 448 0 0 0 io_oeb[1]
port 15 nsew signal tristate
flabel metal2 s 25536 79200 25648 80000 0 FreeSans 448 90 0 0 io_oeb[20]
port 16 nsew signal tristate
flabel metal2 s 30240 79200 30352 80000 0 FreeSans 448 90 0 0 io_oeb[21]
port 17 nsew signal tristate
flabel metal2 s 34272 79200 34384 80000 0 FreeSans 448 90 0 0 io_oeb[22]
port 18 nsew signal tristate
flabel metal2 s 58464 79200 58576 80000 0 FreeSans 448 90 0 0 io_oeb[23]
port 19 nsew signal tristate
flabel metal3 s 79200 57792 80000 57904 0 FreeSans 448 0 0 0 io_oeb[24]
port 20 nsew signal tristate
flabel metal3 s 79200 16128 80000 16240 0 FreeSans 448 0 0 0 io_oeb[25]
port 21 nsew signal tristate
flabel metal3 s 79200 19488 80000 19600 0 FreeSans 448 0 0 0 io_oeb[26]
port 22 nsew signal tristate
flabel metal3 s 79200 64512 80000 64624 0 FreeSans 448 0 0 0 io_oeb[27]
port 23 nsew signal tristate
flabel metal3 s 79200 28224 80000 28336 0 FreeSans 448 0 0 0 io_oeb[28]
port 24 nsew signal tristate
flabel metal3 s 79200 46368 80000 46480 0 FreeSans 448 0 0 0 io_oeb[29]
port 25 nsew signal tristate
flabel metal2 s 56448 79200 56560 80000 0 FreeSans 448 90 0 0 io_oeb[2]
port 26 nsew signal tristate
flabel metal2 s 63168 0 63280 800 0 FreeSans 448 90 0 0 io_oeb[30]
port 27 nsew signal tristate
flabel metal2 s 60480 79200 60592 80000 0 FreeSans 448 90 0 0 io_oeb[31]
port 28 nsew signal tristate
flabel metal3 s 79200 59808 80000 59920 0 FreeSans 448 0 0 0 io_oeb[32]
port 29 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 io_oeb[33]
port 30 nsew signal tristate
flabel metal2 s 59136 0 59248 800 0 FreeSans 448 90 0 0 io_oeb[34]
port 31 nsew signal tristate
flabel metal2 s 49728 79200 49840 80000 0 FreeSans 448 90 0 0 io_oeb[35]
port 32 nsew signal tristate
flabel metal2 s 59808 79200 59920 80000 0 FreeSans 448 90 0 0 io_oeb[36]
port 33 nsew signal tristate
flabel metal2 s 49728 0 49840 800 0 FreeSans 448 90 0 0 io_oeb[37]
port 34 nsew signal tristate
flabel metal2 s 35616 79200 35728 80000 0 FreeSans 448 90 0 0 io_oeb[3]
port 35 nsew signal tristate
flabel metal2 s 34944 79200 35056 80000 0 FreeSans 448 90 0 0 io_oeb[4]
port 36 nsew signal tristate
flabel metal3 s 79200 60480 80000 60592 0 FreeSans 448 0 0 0 io_oeb[5]
port 37 nsew signal tristate
flabel metal3 s 79200 18816 80000 18928 0 FreeSans 448 0 0 0 io_oeb[6]
port 38 nsew signal tristate
flabel metal3 s 79200 15456 80000 15568 0 FreeSans 448 0 0 0 io_oeb[7]
port 39 nsew signal tristate
flabel metal2 s 57792 79200 57904 80000 0 FreeSans 448 90 0 0 io_oeb[8]
port 40 nsew signal tristate
flabel metal3 s 79200 37632 80000 37744 0 FreeSans 448 0 0 0 io_oeb[9]
port 41 nsew signal tristate
flabel metal3 s 79200 40320 80000 40432 0 FreeSans 448 0 0 0 rst
port 42 nsew signal input
flabel metal3 s 79200 42336 80000 42448 0 FreeSans 448 0 0 0 salida[0]
port 43 nsew signal tristate
flabel metal3 s 79200 45024 80000 45136 0 FreeSans 448 0 0 0 salida[1]
port 44 nsew signal tristate
flabel metal2 s 47040 79200 47152 80000 0 FreeSans 448 90 0 0 salida[2]
port 45 nsew signal tristate
flabel metal3 s 79200 47712 80000 47824 0 FreeSans 448 0 0 0 salida[3]
port 46 nsew signal tristate
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 47 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 47 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 47 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 48 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 48 nsew ground bidirectional
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal3 36288 36680 36288 36680 0 _000_
rlabel metal2 34328 37240 34328 37240 0 _001_
rlabel metal2 41272 39088 41272 39088 0 _002_
rlabel metal2 39816 34496 39816 34496 0 _003_
rlabel metal2 43288 36176 43288 36176 0 _004_
rlabel metal2 43176 32200 43176 32200 0 _005_
rlabel metal2 42448 29960 42448 29960 0 _006_
rlabel metal2 37464 32256 37464 32256 0 _007_
rlabel metal2 38304 27944 38304 27944 0 _008_
rlabel metal2 39872 28728 39872 28728 0 _009_
rlabel metal2 34776 28560 34776 28560 0 _010_
rlabel metal2 33432 28952 33432 28952 0 _011_
rlabel metal2 30184 28952 30184 28952 0 _012_
rlabel metal2 33656 32704 33656 32704 0 _013_
rlabel metal2 28840 31304 28840 31304 0 _014_
rlabel metal2 31416 34552 31416 34552 0 _015_
rlabel metal2 29736 37744 29736 37744 0 _016_
rlabel metal2 30352 38920 30352 38920 0 _017_
rlabel metal2 28728 41608 28728 41608 0 _018_
rlabel metal2 29960 43064 29960 43064 0 _019_
rlabel metal2 29176 46984 29176 46984 0 _020_
rlabel metal2 31640 45248 31640 45248 0 _021_
rlabel metal2 34552 47096 34552 47096 0 _022_
rlabel metal2 37632 46088 37632 46088 0 _023_
rlabel metal2 38808 45528 38808 45528 0 _024_
rlabel metal3 40600 41272 40600 41272 0 _025_
rlabel metal2 41048 41160 41048 41160 0 _026_
rlabel metal2 51464 42336 51464 42336 0 _027_
rlabel metal3 51856 45080 51856 45080 0 _028_
rlabel metal2 45640 48664 45640 48664 0 _029_
rlabel metal2 51576 47824 51576 47824 0 _030_
rlabel metal2 43400 44296 43400 44296 0 _031_
rlabel metal3 44800 46536 44800 46536 0 _032_
rlabel metal3 43792 44184 43792 44184 0 _033_
rlabel metal3 48776 40488 48776 40488 0 _034_
rlabel metal2 46536 40432 46536 40432 0 _035_
rlabel metal2 45976 41608 45976 41608 0 _036_
rlabel metal2 43400 40712 43400 40712 0 _037_
rlabel metal3 36288 38696 36288 38696 0 _038_
rlabel metal2 35448 39200 35448 39200 0 _039_
rlabel metal2 34664 46984 34664 46984 0 _040_
rlabel metal2 40040 37240 40040 37240 0 _041_
rlabel metal2 40656 38808 40656 38808 0 _042_
rlabel metal3 42672 30408 42672 30408 0 _043_
rlabel metal2 41272 34888 41272 34888 0 _044_
rlabel metal2 40152 33600 40152 33600 0 _045_
rlabel metal2 40264 35168 40264 35168 0 _046_
rlabel metal2 42952 35728 42952 35728 0 _047_
rlabel metal2 42000 31752 42000 31752 0 _048_
rlabel metal2 45080 32592 45080 32592 0 _049_
rlabel metal2 43400 32984 43400 32984 0 _050_
rlabel metal2 42280 30240 42280 30240 0 _051_
rlabel metal2 42336 30408 42336 30408 0 _052_
rlabel metal2 37576 31360 37576 31360 0 _053_
rlabel metal2 37800 31696 37800 31696 0 _054_
rlabel metal2 38584 31808 38584 31808 0 _055_
rlabel metal2 38696 28952 38696 28952 0 _056_
rlabel metal3 40320 28056 40320 28056 0 _057_
rlabel metal2 40040 29904 40040 29904 0 _058_
rlabel metal2 37800 28224 37800 28224 0 _059_
rlabel metal3 34384 29400 34384 29400 0 _060_
rlabel metal2 37128 27216 37128 27216 0 _061_
rlabel metal2 36176 28840 36176 28840 0 _062_
rlabel metal2 36232 30296 36232 30296 0 _063_
rlabel metal3 35784 31192 35784 31192 0 _064_
rlabel metal3 32984 29176 32984 29176 0 _065_
rlabel metal2 36008 28784 36008 28784 0 _066_
rlabel metal2 31528 28448 31528 28448 0 _067_
rlabel metal2 32424 31752 32424 31752 0 _068_
rlabel metal2 32592 32312 32592 32312 0 _069_
rlabel metal2 31304 33376 31304 33376 0 _070_
rlabel metal2 30744 32144 30744 32144 0 _071_
rlabel metal2 32928 33544 32928 33544 0 _072_
rlabel metal2 31640 39984 31640 39984 0 _073_
rlabel metal2 31416 33656 31416 33656 0 _074_
rlabel metal2 30576 37912 30576 37912 0 _075_
rlabel metal2 30744 40712 30744 40712 0 _076_
rlabel metal2 30632 39872 30632 39872 0 _077_
rlabel metal2 32088 39928 32088 39928 0 _078_
rlabel metal3 31808 41720 31808 41720 0 _079_
rlabel metal2 31192 42728 31192 42728 0 _080_
rlabel metal2 31192 41272 31192 41272 0 _081_
rlabel metal2 33992 43456 33992 43456 0 _082_
rlabel metal2 30968 45864 30968 45864 0 _083_
rlabel metal2 31528 43512 31528 43512 0 _084_
rlabel metal2 30632 46088 30632 46088 0 _085_
rlabel metal2 31920 45080 31920 45080 0 _086_
rlabel metal2 34440 45584 34440 45584 0 _087_
rlabel metal2 33208 46088 33208 46088 0 _088_
rlabel metal2 34272 46536 34272 46536 0 _089_
rlabel metal2 39256 44576 39256 44576 0 _090_
rlabel metal2 35448 45752 35448 45752 0 _091_
rlabel metal2 39928 43904 39928 43904 0 _092_
rlabel metal2 37912 44184 37912 44184 0 _093_
rlabel metal2 39816 44632 39816 44632 0 _094_
rlabel metal2 39144 45080 39144 45080 0 _095_
rlabel metal2 38136 42336 38136 42336 0 _096_
rlabel metal3 39088 41384 39088 41384 0 _097_
rlabel metal2 39368 43568 39368 43568 0 _098_
rlabel metal3 41160 41888 41160 41888 0 _099_
rlabel metal2 38360 42224 38360 42224 0 _100_
rlabel metal2 51464 44072 51464 44072 0 _101_
rlabel metal2 51912 47096 51912 47096 0 _102_
rlabel metal2 50904 46312 50904 46312 0 _103_
rlabel metal2 51688 45584 51688 45584 0 _104_
rlabel metal2 50456 44408 50456 44408 0 _105_
rlabel metal2 47656 46144 47656 46144 0 _106_
rlabel metal2 50232 47488 50232 47488 0 _107_
rlabel metal2 47880 47264 47880 47264 0 _108_
rlabel metal2 52696 44912 52696 44912 0 _109_
rlabel metal3 52360 42952 52360 42952 0 _110_
rlabel metal2 50344 45136 50344 45136 0 _111_
rlabel metal2 52976 44072 52976 44072 0 _112_
rlabel metal3 45696 45192 45696 45192 0 _113_
rlabel metal2 46424 47824 46424 47824 0 _114_
rlabel metal3 52248 47320 52248 47320 0 _115_
rlabel metal3 51296 46872 51296 46872 0 _116_
rlabel metal3 46480 45080 46480 45080 0 _117_
rlabel metal2 46424 44800 46424 44800 0 _118_
rlabel metal2 45640 47152 45640 47152 0 _119_
rlabel metal3 48216 48440 48216 48440 0 _120_
rlabel metal2 47432 46088 47432 46088 0 _121_
rlabel metal2 48440 45864 48440 45864 0 _122_
rlabel metal2 46704 46872 46704 46872 0 _123_
rlabel metal2 48440 46256 48440 46256 0 _124_
rlabel metal2 49224 47712 49224 47712 0 _125_
rlabel metal2 48328 47320 48328 47320 0 _126_
rlabel metal2 46872 47040 46872 47040 0 _127_
rlabel metal2 45696 44184 45696 44184 0 _128_
rlabel metal3 48720 46760 48720 46760 0 _129_
rlabel metal3 48496 46088 48496 46088 0 _130_
rlabel metal2 45864 44520 45864 44520 0 _131_
rlabel metal2 45864 41160 45864 41160 0 _132_
rlabel metal2 47768 41440 47768 41440 0 _133_
rlabel metal2 43624 40432 43624 40432 0 _134_
rlabel metal2 37968 39032 37968 39032 0 _135_
rlabel metal2 33712 45080 33712 45080 0 _136_
rlabel metal2 33320 44016 33320 44016 0 _137_
rlabel metal2 33096 41160 33096 41160 0 _138_
rlabel metal2 38920 42224 38920 42224 0 _139_
rlabel metal2 39480 37352 39480 37352 0 _140_
rlabel metal2 39592 36960 39592 36960 0 _141_
rlabel metal2 39592 29624 39592 29624 0 _142_
rlabel metal2 39704 37128 39704 37128 0 _143_
rlabel metal2 32536 34440 32536 34440 0 _144_
rlabel metal2 32424 33600 32424 33600 0 _145_
rlabel metal2 38472 30856 38472 30856 0 _146_
rlabel metal2 35896 31416 35896 31416 0 _147_
rlabel metal2 35728 33208 35728 33208 0 _148_
rlabel metal2 40040 33824 40040 33824 0 _149_
rlabel metal2 40376 38024 40376 38024 0 _150_
rlabel metal2 41720 40824 41720 40824 0 _151_
rlabel metal2 39816 43568 39816 43568 0 _152_
rlabel metal2 42616 36344 42616 36344 0 _153_
rlabel metal2 28280 2478 28280 2478 0 clk
rlabel metal2 77336 40712 77336 40712 0 clk_s
rlabel metal2 39256 35728 39256 35728 0 clknet_0_clk
rlabel metal2 29176 36064 29176 36064 0 clknet_2_0__leaf_clk
rlabel metal2 39144 29792 39144 29792 0 clknet_2_1__leaf_clk
rlabel metal2 29288 42280 29288 42280 0 clknet_2_2__leaf_clk
rlabel metal2 42168 46648 42168 46648 0 clknet_2_3__leaf_clk
rlabel metal2 38024 38724 38024 38724 0 count\[0\]
rlabel metal2 36960 27720 36960 27720 0 count\[10\]
rlabel metal2 36120 30352 36120 30352 0 count\[11\]
rlabel metal2 31976 32760 31976 32760 0 count\[12\]
rlabel metal2 32200 32704 32200 32704 0 count\[13\]
rlabel metal2 30968 31696 30968 31696 0 count\[14\]
rlabel metal2 32312 33152 32312 33152 0 count\[15\]
rlabel metal2 32648 39536 32648 39536 0 count\[16\]
rlabel metal2 32424 40096 32424 40096 0 count\[17\]
rlabel metal3 33096 41944 33096 41944 0 count\[18\]
rlabel metal2 32088 43176 32088 43176 0 count\[19\]
rlabel metal2 39144 36624 39144 36624 0 count\[1\]
rlabel metal2 31304 45808 31304 45808 0 count\[20\]
rlabel metal2 33376 45864 33376 45864 0 count\[21\]
rlabel metal2 34664 44744 34664 44744 0 count\[22\]
rlabel metal2 34776 44576 34776 44576 0 count\[23\]
rlabel metal2 39592 45192 39592 45192 0 count\[24\]
rlabel metal2 38696 43848 38696 43848 0 count\[25\]
rlabel metal2 39144 42000 39144 42000 0 count\[26\]
rlabel metal2 40376 36400 40376 36400 0 count\[2\]
rlabel metal2 41440 36456 41440 36456 0 count\[3\]
rlabel metal2 42280 35672 42280 35672 0 count\[4\]
rlabel metal2 42168 34160 42168 34160 0 count\[5\]
rlabel metal2 44856 31304 44856 31304 0 count\[6\]
rlabel metal2 39368 31752 39368 31752 0 count\[7\]
rlabel metal2 39816 29512 39816 29512 0 count\[8\]
rlabel via2 41048 28728 41048 28728 0 count\[9\]
rlabel metal2 78232 47152 78232 47152 0 dir
rlabel metal3 78722 45752 78722 45752 0 enable
rlabel metal2 50568 47880 50568 47880 0 net1
rlabel metal2 51464 45304 51464 45304 0 net10
rlabel metal2 45640 42224 45640 42224 0 net11
rlabel metal2 75656 40488 75656 40488 0 net12
rlabel metal2 78232 15680 78232 15680 0 net13
rlabel metal2 57960 76664 57960 76664 0 net14
rlabel metal2 78232 37744 78232 37744 0 net15
rlabel metal2 48440 2030 48440 2030 0 net16
rlabel metal2 62552 2030 62552 2030 0 net17
rlabel metal2 78232 50064 78232 50064 0 net18
rlabel metal2 59304 76664 59304 76664 0 net19
rlabel metal2 50512 47208 50512 47208 0 net2
rlabel metal2 51240 76944 51240 76944 0 net20
rlabel metal2 78232 29232 78232 29232 0 net21
rlabel metal2 67256 2030 67256 2030 0 net22
rlabel metal2 78288 17416 78288 17416 0 net23
rlabel metal2 38360 2030 38360 2030 0 net24
rlabel metal3 78736 43736 78736 43736 0 net25
rlabel metal2 25704 76664 25704 76664 0 net26
rlabel metal2 30408 76664 30408 76664 0 net27
rlabel metal2 34440 76664 34440 76664 0 net28
rlabel metal2 58688 76664 58688 76664 0 net29
rlabel metal2 77896 41104 77896 41104 0 net3
rlabel metal2 78232 58016 78232 58016 0 net30
rlabel metal2 78232 16576 78232 16576 0 net31
rlabel metal3 78736 20216 78736 20216 0 net32
rlabel metal3 78722 64568 78722 64568 0 net33
rlabel metal2 78232 28336 78232 28336 0 net34
rlabel metal2 78232 46592 78232 46592 0 net35
rlabel metal2 63224 2030 63224 2030 0 net36
rlabel metal2 60648 76664 60648 76664 0 net37
rlabel metal3 78722 59864 78722 59864 0 net38
rlabel metal2 35000 2030 35000 2030 0 net39
rlabel metal2 45528 40488 45528 40488 0 net4
rlabel metal2 59192 2030 59192 2030 0 net40
rlabel metal2 50344 76832 50344 76832 0 net41
rlabel metal2 59976 76664 59976 76664 0 net42
rlabel metal2 49784 2030 49784 2030 0 net43
rlabel metal2 78232 27048 78232 27048 0 net44
rlabel metal2 78232 30016 78232 30016 0 net45
rlabel metal2 56616 76328 56616 76328 0 net46
rlabel metal2 36008 77000 36008 77000 0 net47
rlabel metal2 35112 76328 35112 76328 0 net48
rlabel metal3 78722 60536 78722 60536 0 net49
rlabel metal2 53536 42504 53536 42504 0 net5
rlabel metal2 78232 19096 78232 19096 0 net50
rlabel metal2 53368 44688 53368 44688 0 net6
rlabel metal2 50120 76440 50120 76440 0 net7
rlabel metal2 52808 47376 52808 47376 0 net8
rlabel metal2 45248 41944 45248 41944 0 net9
rlabel metal2 78232 40712 78232 40712 0 rst
rlabel metal2 78008 42112 78008 42112 0 salida[0]
rlabel metal2 78008 45024 78008 45024 0 salida[1]
rlabel metal2 47096 77770 47096 77770 0 salida[2]
rlabel metal2 78008 47880 78008 47880 0 salida[3]
rlabel metal2 50792 42616 50792 42616 0 state\[0\]
rlabel metal2 51688 42560 51688 42560 0 state\[1\]
rlabel metal2 51296 43736 51296 43736 0 state\[2\]
rlabel metal2 46424 43512 46424 43512 0 state_next\[0\]
rlabel metal2 45192 46928 45192 46928 0 state_next\[1\]
rlabel metal2 44576 44408 44576 44408 0 state_next\[2\]
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
