module control_system (clk,
    clk_s,
    dir,
    enable,
    rst,
    vdd,
    vss,
    io_oeb,
    salida);
 input clk;
 output clk_s;
 input dir;
 input enable;
 input rst;
 input vdd;
 input vss;
 output [37:0] io_oeb;
 output [3:0] salida;

 wire net44;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net45;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net46;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net13;
 wire net14;
 wire net15;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire \count[0] ;
 wire \count[10] ;
 wire \count[11] ;
 wire \count[12] ;
 wire \count[13] ;
 wire \count[14] ;
 wire \count[15] ;
 wire \count[16] ;
 wire \count[17] ;
 wire \count[18] ;
 wire \count[19] ;
 wire \count[1] ;
 wire \count[20] ;
 wire \count[21] ;
 wire \count[22] ;
 wire \count[23] ;
 wire \count[24] ;
 wire \count[25] ;
 wire \count[26] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \count[5] ;
 wire \count[6] ;
 wire \count[7] ;
 wire \count[8] ;
 wire \count[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state_next[0] ;
 wire \state_next[1] ;
 wire \state_next[2] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__A1 (.I(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A1 (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A1 (.I(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A1 (.I(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__I (.I(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__A1 (.I(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__I (.I(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__A1 (.I(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__A2 (.I(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__A1 (.I(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__I (.I(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A2 (.I(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__I (.I(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout11_I (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(dir),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(enable),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(rst),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output4_I (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output5_I (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_420 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_425 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_537 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_541 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_573 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_588 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_611 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_446 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_675 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_468 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_462 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_320 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_480 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_421 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_429 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_462 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_474 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_675 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_677 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_446 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_497 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_513 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_675 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_490 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_497 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_509 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_533 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_541 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _154_ (.I(\count[0] ),
    .Z(_135_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _155_ (.I(\count[22] ),
    .ZN(_136_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _156_ (.A1(\count[20] ),
    .A2(\count[21] ),
    .A3(_136_),
    .A4(\count[23] ),
    .ZN(_137_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _157_ (.A1(\count[16] ),
    .A2(\count[17] ),
    .ZN(_138_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _158_ (.A1(\count[18] ),
    .A2(\count[19] ),
    .A3(_137_),
    .A4(_138_),
    .ZN(_139_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _159_ (.A1(\count[24] ),
    .A2(\count[25] ),
    .A3(\count[26] ),
    .A4(_139_),
    .ZN(_140_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _160_ (.A1(\count[2] ),
    .A2(\count[3] ),
    .A3(\count[4] ),
    .A4(\count[5] ),
    .ZN(_141_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _161_ (.A1(\count[8] ),
    .A2(\count[9] ),
    .ZN(_142_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _162_ (.A1(_135_),
    .A2(\count[1] ),
    .A3(_142_),
    .ZN(_143_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _163_ (.I(\count[15] ),
    .ZN(_144_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _164_ (.A1(\count[14] ),
    .A2(_144_),
    .ZN(_145_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _165_ (.I(\count[7] ),
    .ZN(_146_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _166_ (.I(\count[10] ),
    .ZN(_147_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _167_ (.A1(\count[6] ),
    .A2(_146_),
    .A3(_147_),
    .A4(\count[11] ),
    .ZN(_148_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _168_ (.A1(\count[12] ),
    .A2(\count[13] ),
    .A3(_145_),
    .A4(_148_),
    .ZN(_149_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _169_ (.A1(_140_),
    .A2(_141_),
    .A3(_143_),
    .A4(_149_),
    .Z(_150_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _170_ (.A1(net3),
    .A2(_150_),
    .Z(_151_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _171_ (.I(_151_),
    .Z(_152_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _172_ (.I(_152_),
    .Z(_153_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _173_ (.A1(_135_),
    .A2(_153_),
    .ZN(_000_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _174_ (.A1(_135_),
    .A2(\count[1] ),
    .ZN(_038_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _175_ (.I(_151_),
    .Z(_039_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _176_ (.I(_039_),
    .Z(_040_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _177_ (.A1(_135_),
    .A2(\count[1] ),
    .Z(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _178_ (.A1(_038_),
    .A2(_040_),
    .A3(_041_),
    .ZN(_001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _179_ (.A1(\count[2] ),
    .A2(_041_),
    .ZN(_042_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _180_ (.A1(_153_),
    .A2(_042_),
    .ZN(_002_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _181_ (.I(_039_),
    .Z(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _182_ (.A1(\count[0] ),
    .A2(\count[1] ),
    .A3(\count[2] ),
    .A4(\count[3] ),
    .Z(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _183_ (.I(_044_),
    .Z(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _184_ (.A1(\count[2] ),
    .A2(_041_),
    .B(\count[3] ),
    .ZN(_046_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _185_ (.A1(_043_),
    .A2(_045_),
    .A3(_046_),
    .ZN(_003_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _186_ (.A1(\count[4] ),
    .A2(_045_),
    .ZN(_047_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _187_ (.A1(_153_),
    .A2(_047_),
    .ZN(_004_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _188_ (.A1(\count[4] ),
    .A2(\count[5] ),
    .Z(_048_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _189_ (.A1(_045_),
    .A2(_048_),
    .Z(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _190_ (.A1(\count[4] ),
    .A2(_045_),
    .B(\count[5] ),
    .ZN(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _191_ (.A1(_043_),
    .A2(_049_),
    .A3(_050_),
    .ZN(_005_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _192_ (.A1(\count[6] ),
    .A2(_049_),
    .Z(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _193_ (.A1(\count[6] ),
    .A2(_049_),
    .ZN(_052_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _194_ (.A1(_043_),
    .A2(_051_),
    .A3(_052_),
    .ZN(_006_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _195_ (.I(_039_),
    .Z(_053_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _196_ (.A1(_146_),
    .A2(_051_),
    .Z(_054_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _197_ (.A1(_053_),
    .A2(_054_),
    .ZN(_007_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _198_ (.A1(\count[6] ),
    .A2(\count[7] ),
    .A3(_044_),
    .A4(_048_),
    .ZN(_055_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _199_ (.A1(\count[8] ),
    .A2(_055_),
    .Z(_056_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _200_ (.A1(_053_),
    .A2(_056_),
    .ZN(_008_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _201_ (.I(\count[9] ),
    .ZN(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _202_ (.A1(\count[7] ),
    .A2(\count[8] ),
    .A3(_051_),
    .ZN(_058_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _203_ (.A1(_142_),
    .A2(_055_),
    .ZN(_059_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _204_ (.A1(_057_),
    .A2(_058_),
    .B(_059_),
    .C(_043_),
    .ZN(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _205_ (.I(_039_),
    .Z(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _206_ (.A1(\count[10] ),
    .A2(_059_),
    .ZN(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _207_ (.A1(_147_),
    .A2(_142_),
    .A3(_055_),
    .ZN(_062_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _208_ (.A1(_060_),
    .A2(_061_),
    .A3(_062_),
    .ZN(_010_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _209_ (.I(\count[11] ),
    .ZN(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _210_ (.A1(_147_),
    .A2(_063_),
    .A3(_142_),
    .A4(_055_),
    .ZN(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _211_ (.I(_064_),
    .Z(_065_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _212_ (.A1(\count[11] ),
    .A2(_062_),
    .ZN(_066_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _213_ (.A1(_060_),
    .A2(_065_),
    .A3(_066_),
    .ZN(_011_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _214_ (.A1(\count[12] ),
    .A2(_065_),
    .ZN(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _215_ (.A1(_053_),
    .A2(_067_),
    .ZN(_012_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _216_ (.A1(\count[12] ),
    .A2(_065_),
    .B(\count[13] ),
    .ZN(_068_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _217_ (.A1(\count[12] ),
    .A2(\count[13] ),
    .Z(_069_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _218_ (.A1(_065_),
    .A2(_069_),
    .Z(_070_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _219_ (.A1(_060_),
    .A2(_068_),
    .A3(_070_),
    .ZN(_013_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _220_ (.A1(\count[14] ),
    .A2(_070_),
    .ZN(_071_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _221_ (.A1(_053_),
    .A2(_071_),
    .ZN(_014_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _222_ (.A1(\count[14] ),
    .A2(\count[15] ),
    .A3(_064_),
    .A4(_069_),
    .Z(_072_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _223_ (.I(_072_),
    .Z(_073_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _224_ (.A1(\count[14] ),
    .A2(_070_),
    .B(\count[15] ),
    .ZN(_074_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _225_ (.A1(_060_),
    .A2(_073_),
    .A3(_074_),
    .ZN(_015_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _226_ (.A1(\count[16] ),
    .A2(_073_),
    .ZN(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _227_ (.A1(_040_),
    .A2(_075_),
    .ZN(_016_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _228_ (.I(_151_),
    .Z(_076_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _229_ (.A1(\count[16] ),
    .A2(_073_),
    .B(\count[17] ),
    .ZN(_077_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _230_ (.A1(\count[16] ),
    .A2(\count[17] ),
    .Z(_078_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _231_ (.A1(_073_),
    .A2(_078_),
    .Z(_079_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _232_ (.A1(_076_),
    .A2(_077_),
    .A3(_079_),
    .ZN(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _233_ (.A1(\count[18] ),
    .A2(_079_),
    .Z(_080_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _234_ (.A1(\count[18] ),
    .A2(_079_),
    .ZN(_081_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _235_ (.A1(_076_),
    .A2(_080_),
    .A3(_081_),
    .ZN(_018_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _236_ (.A1(\count[18] ),
    .A2(\count[19] ),
    .A3(_072_),
    .A4(_078_),
    .Z(_082_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _237_ (.I(_082_),
    .Z(_083_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _238_ (.A1(\count[19] ),
    .A2(_080_),
    .ZN(_084_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _239_ (.A1(_076_),
    .A2(_083_),
    .A3(_084_),
    .ZN(_019_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _240_ (.A1(\count[20] ),
    .A2(_083_),
    .ZN(_085_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _241_ (.A1(_040_),
    .A2(_085_),
    .ZN(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _242_ (.A1(\count[20] ),
    .A2(_083_),
    .B(\count[21] ),
    .ZN(_086_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _243_ (.A1(\count[20] ),
    .A2(\count[21] ),
    .Z(_087_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _244_ (.A1(_082_),
    .A2(_087_),
    .Z(_088_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _245_ (.A1(_076_),
    .A2(_086_),
    .A3(_088_),
    .ZN(_021_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _246_ (.A1(_136_),
    .A2(_088_),
    .Z(_089_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _247_ (.A1(_040_),
    .A2(_089_),
    .ZN(_022_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _248_ (.A1(\count[22] ),
    .A2(\count[23] ),
    .A3(_083_),
    .A4(_087_),
    .Z(_090_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _249_ (.A1(\count[22] ),
    .A2(_088_),
    .B(\count[23] ),
    .ZN(_091_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _250_ (.A1(_152_),
    .A2(_090_),
    .A3(_091_),
    .ZN(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _251_ (.I(\count[24] ),
    .ZN(_092_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _252_ (.A1(\count[22] ),
    .A2(\count[23] ),
    .A3(_082_),
    .A4(_087_),
    .ZN(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _253_ (.A1(_092_),
    .A2(_093_),
    .ZN(_094_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _254_ (.A1(\count[24] ),
    .A2(_090_),
    .ZN(_095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _255_ (.A1(_152_),
    .A2(_094_),
    .A3(_095_),
    .ZN(_024_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _256_ (.I(\count[25] ),
    .ZN(_096_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _257_ (.A1(_092_),
    .A2(_096_),
    .A3(_093_),
    .ZN(_097_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _258_ (.A1(\count[24] ),
    .A2(_090_),
    .B(\count[25] ),
    .ZN(_098_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _259_ (.A1(_152_),
    .A2(_097_),
    .A3(_098_),
    .ZN(_025_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _260_ (.A1(_092_),
    .A2(_096_),
    .A3(_093_),
    .B(\count[26] ),
    .ZN(_099_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _261_ (.A1(_092_),
    .A2(_096_),
    .A3(\count[26] ),
    .A4(_093_),
    .Z(_100_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _262_ (.A1(_099_),
    .A2(_100_),
    .B(_153_),
    .ZN(_026_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _263_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .ZN(_101_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _264_ (.A1(\state[2] ),
    .A2(_101_),
    .ZN(_102_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _265_ (.A1(\state[2] ),
    .A2(_101_),
    .ZN(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _266_ (.I(\state[0] ),
    .Z(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _267_ (.I(\state[2] ),
    .ZN(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _268_ (.A1(\state[1] ),
    .A2(_104_),
    .A3(_105_),
    .ZN(_106_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _269_ (.A1(_103_),
    .A2(_106_),
    .ZN(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _270_ (.A1(_102_),
    .A2(_107_),
    .ZN(_108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _271_ (.I(_108_),
    .Z(_109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _272_ (.A1(net5),
    .A2(_109_),
    .ZN(_110_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _273_ (.A1(\state[1] ),
    .A2(\state[2] ),
    .A3(_101_),
    .B(_110_),
    .ZN(_027_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _274_ (.A1(\state[1] ),
    .A2(_105_),
    .ZN(_111_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _275_ (.A1(net6),
    .A2(_109_),
    .ZN(_112_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _276_ (.A1(_104_),
    .A2(_111_),
    .B(_112_),
    .ZN(_028_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _277_ (.I(_108_),
    .Z(_113_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _278_ (.A1(net7),
    .A2(_113_),
    .ZN(_114_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _279_ (.A1(_106_),
    .A2(_114_),
    .ZN(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _280_ (.I(net8),
    .ZN(_115_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _281_ (.I(_103_),
    .Z(_116_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _282_ (.A1(_115_),
    .A2(_116_),
    .B(_102_),
    .ZN(_030_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _283_ (.A1(net2),
    .A2(_104_),
    .ZN(_117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _284_ (.A1(\state_next[0] ),
    .A2(_109_),
    .ZN(_118_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _285_ (.A1(_113_),
    .A2(_117_),
    .B(_118_),
    .ZN(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _286_ (.I(\state_next[1] ),
    .ZN(_119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _287_ (.I(net2),
    .Z(_120_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _288_ (.I(_106_),
    .ZN(_121_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _289_ (.A1(net1),
    .A2(net2),
    .ZN(_122_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _290_ (.A1(_120_),
    .A2(_121_),
    .B(_107_),
    .C(_122_),
    .ZN(_123_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _291_ (.A1(net1),
    .A2(_120_),
    .A3(_116_),
    .A4(_111_),
    .Z(_124_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _292_ (.I(net1),
    .ZN(_125_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _293_ (.A1(_125_),
    .A2(_120_),
    .B(_104_),
    .C(_111_),
    .ZN(_126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _294_ (.A1(_108_),
    .A2(_124_),
    .A3(_126_),
    .ZN(_127_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _295_ (.A1(_119_),
    .A2(_113_),
    .B1(_123_),
    .B2(_127_),
    .ZN(_032_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _296_ (.I(\state_next[2] ),
    .ZN(_128_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _297_ (.A1(_125_),
    .A2(net2),
    .A3(_116_),
    .A4(_111_),
    .ZN(_129_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _298_ (.A1(_120_),
    .A2(_116_),
    .B1(_106_),
    .B2(_122_),
    .C(_129_),
    .ZN(_130_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _299_ (.A1(_109_),
    .A2(_130_),
    .ZN(_131_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _300_ (.A1(_128_),
    .A2(_113_),
    .B(_131_),
    .ZN(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _301_ (.I(net3),
    .Z(_132_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _302_ (.A1(_132_),
    .A2(\state_next[0] ),
    .Z(_133_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _303_ (.I(_133_),
    .Z(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _304_ (.A1(_132_),
    .A2(_119_),
    .ZN(_035_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _305_ (.A1(_132_),
    .A2(_128_),
    .ZN(_036_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _306_ (.A1(net9),
    .A2(_150_),
    .ZN(_134_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _307_ (.A1(_132_),
    .A2(_134_),
    .ZN(_037_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _308_ (.D(_000_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _309_ (.D(_001_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _310_ (.D(_002_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _311_ (.D(_003_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _312_ (.D(_004_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _313_ (.D(_005_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _314_ (.D(_006_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _315_ (.D(_007_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _316_ (.D(_008_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _317_ (.D(_009_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _318_ (.D(_010_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _319_ (.D(_011_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _320_ (.D(_012_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[12] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _321_ (.D(_013_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[13] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _322_ (.D(_014_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[14] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _323_ (.D(_015_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[15] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _324_ (.D(_016_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[16] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _325_ (.D(_017_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[17] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _326_ (.D(_018_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[18] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _327_ (.D(_019_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[19] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _328_ (.D(_020_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[20] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _329_ (.D(_021_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[21] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _330_ (.D(_022_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[22] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _331_ (.D(_023_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[23] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _332_ (.D(_024_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[24] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _333_ (.D(_025_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[25] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _334_ (.D(_026_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[26] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _335_ (.D(_027_),
    .CLK(net10),
    .Q(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _336_ (.D(_028_),
    .CLK(net10),
    .Q(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _337_ (.D(_029_),
    .CLK(net9),
    .Q(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _338_ (.D(_030_),
    .CLK(net10),
    .Q(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _339_ (.D(_031_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state_next[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _340_ (.D(_032_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state_next[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _341_ (.D(_033_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state_next[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _342_ (.D(_034_),
    .CLK(net10),
    .Q(\state[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _343_ (.D(_035_),
    .CLK(net9),
    .Q(\state[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _344_ (.D(_036_),
    .CLK(net9),
    .Q(\state[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _345_ (.D(_037_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_13 (.ZN(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_14 (.ZN(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_15 (.ZN(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_16 (.ZN(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_17 (.ZN(net17),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_18 (.ZN(net18),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_19 (.ZN(net19),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_20 (.ZN(net20),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_21 (.ZN(net21),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_22 (.ZN(net22),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_23 (.ZN(net23),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_24 (.ZN(net24),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_25 (.ZN(net25),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_26 (.ZN(net26),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_27 (.ZN(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_28 (.ZN(net28),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_29 (.ZN(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_30 (.ZN(net30),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_31 (.ZN(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_32 (.ZN(net32),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_33 (.ZN(net33),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_34 (.ZN(net34),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_35 (.ZN(net35),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_36 (.ZN(net36),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_37 (.ZN(net37),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_38 (.ZN(net38),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_39 (.ZN(net39),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_40 (.ZN(net40),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_41 (.ZN(net41),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_42 (.ZN(net42),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_43 (.ZN(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_44 (.Z(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_45 (.Z(net45),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_46 (.Z(net46),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_47 (.Z(net47),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_48 (.Z(net48),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_49 (.Z(net49),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_50 (.Z(net50),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout10 (.I(net11),
    .Z(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout11 (.I(net12),
    .Z(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout12 (.I(net4),
    .Z(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout9 (.I(net11),
    .Z(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(dir),
    .Z(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(enable),
    .Z(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(rst),
    .Z(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output4 (.I(net12),
    .Z(clk_s),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output5 (.I(net5),
    .Z(salida[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output6 (.I(net6),
    .Z(salida[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output7 (.I(net7),
    .Z(salida[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output8 (.I(net8),
    .Z(salida[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 assign io_oeb[0] = net44;
 assign io_oeb[10] = net16;
 assign io_oeb[11] = net17;
 assign io_oeb[12] = net18;
 assign io_oeb[13] = net19;
 assign io_oeb[14] = net20;
 assign io_oeb[15] = net21;
 assign io_oeb[16] = net22;
 assign io_oeb[17] = net23;
 assign io_oeb[18] = net24;
 assign io_oeb[19] = net25;
 assign io_oeb[1] = net45;
 assign io_oeb[20] = net26;
 assign io_oeb[21] = net27;
 assign io_oeb[22] = net28;
 assign io_oeb[23] = net29;
 assign io_oeb[24] = net30;
 assign io_oeb[25] = net31;
 assign io_oeb[26] = net32;
 assign io_oeb[27] = net33;
 assign io_oeb[28] = net34;
 assign io_oeb[29] = net35;
 assign io_oeb[2] = net46;
 assign io_oeb[30] = net36;
 assign io_oeb[31] = net37;
 assign io_oeb[32] = net38;
 assign io_oeb[33] = net39;
 assign io_oeb[34] = net40;
 assign io_oeb[35] = net41;
 assign io_oeb[36] = net42;
 assign io_oeb[37] = net43;
 assign io_oeb[3] = net47;
 assign io_oeb[4] = net48;
 assign io_oeb[5] = net49;
 assign io_oeb[6] = net50;
 assign io_oeb[7] = net13;
 assign io_oeb[8] = net14;
 assign io_oeb[9] = net15;
endmodule
