magic
tech gf180mcuD
magscale 1 10
timestamp 1702138370
<< nwell >>
rect 1258 75616 78710 76480
rect 1258 74048 78710 74912
rect 1258 72480 78710 73344
rect 1258 70912 78710 71776
rect 1258 69344 78710 70208
rect 1258 67776 78710 68640
rect 1258 66208 78710 67072
rect 1258 64640 78710 65504
rect 1258 63072 78710 63936
rect 1258 61504 78710 62368
rect 1258 59936 78710 60800
rect 1258 58368 78710 59232
rect 1258 56800 78710 57664
rect 1258 55232 78710 56096
rect 1258 53664 78710 54528
rect 1258 52096 78710 52960
rect 1258 50528 78710 51392
rect 1258 48985 78710 49824
rect 1258 48960 45661 48985
rect 1258 48231 51597 48256
rect 1258 47417 78710 48231
rect 1258 47392 33789 47417
rect 1258 46663 29197 46688
rect 1258 45849 78710 46663
rect 1258 45824 29981 45849
rect 1258 45095 30326 45120
rect 1258 44281 78710 45095
rect 1258 44256 42189 44281
rect 1258 43527 38176 43552
rect 1258 42713 78710 43527
rect 1258 42688 29981 42713
rect 1258 41959 28749 41984
rect 1258 41145 78710 41959
rect 1258 41120 41000 41145
rect 1258 40391 36856 40416
rect 1258 39577 78710 40391
rect 1258 39552 41224 39577
rect 1258 38823 30429 38848
rect 1258 38009 78710 38823
rect 1258 37984 30886 38009
rect 1258 37255 29757 37280
rect 1258 36441 78710 37255
rect 1258 36416 34349 36441
rect 1258 35687 43309 35712
rect 1258 34873 78710 35687
rect 1258 34848 29981 34873
rect 1258 33280 78710 34144
rect 1258 32551 30326 32576
rect 1258 31737 78710 32551
rect 1258 31712 33384 31737
rect 1258 30983 28861 31008
rect 1258 30144 78710 30983
rect 1258 28601 78710 29440
rect 1258 28576 30205 28601
rect 1258 27847 31558 27872
rect 1258 27008 78710 27847
rect 1258 25440 78710 26304
rect 1258 23872 78710 24736
rect 1258 22304 78710 23168
rect 1258 20736 78710 21600
rect 1258 19168 78710 20032
rect 1258 17600 78710 18464
rect 1258 16032 78710 16896
rect 1258 14464 78710 15328
rect 1258 12896 78710 13760
rect 1258 11328 78710 12192
rect 1258 9760 78710 10624
rect 1258 8192 78710 9056
rect 1258 6624 78710 7488
rect 1258 5056 78710 5920
rect 1258 3488 78710 4352
<< pwell >>
rect 1258 76480 78710 76918
rect 1258 74912 78710 75616
rect 1258 73344 78710 74048
rect 1258 71776 78710 72480
rect 1258 70208 78710 70912
rect 1258 68640 78710 69344
rect 1258 67072 78710 67776
rect 1258 65504 78710 66208
rect 1258 63936 78710 64640
rect 1258 62368 78710 63072
rect 1258 60800 78710 61504
rect 1258 59232 78710 59936
rect 1258 57664 78710 58368
rect 1258 56096 78710 56800
rect 1258 54528 78710 55232
rect 1258 52960 78710 53664
rect 1258 51392 78710 52096
rect 1258 49824 78710 50528
rect 1258 48256 78710 48960
rect 1258 46688 78710 47392
rect 1258 45120 78710 45824
rect 1258 43552 78710 44256
rect 1258 41984 78710 42688
rect 1258 40416 78710 41120
rect 1258 38848 78710 39552
rect 1258 37280 78710 37984
rect 1258 35712 78710 36416
rect 1258 34144 78710 34848
rect 1258 32576 78710 33280
rect 1258 31008 78710 31712
rect 1258 29440 78710 30144
rect 1258 27872 78710 28576
rect 1258 26304 78710 27008
rect 1258 24736 78710 25440
rect 1258 23168 78710 23872
rect 1258 21600 78710 22304
rect 1258 20032 78710 20736
rect 1258 18464 78710 19168
rect 1258 16896 78710 17600
rect 1258 15328 78710 16032
rect 1258 13760 78710 14464
rect 1258 12192 78710 12896
rect 1258 10624 78710 11328
rect 1258 9056 78710 9760
rect 1258 7488 78710 8192
rect 1258 5920 78710 6624
rect 1258 4352 78710 5056
rect 1258 3050 78710 3488
<< obsm1 >>
rect 1344 3076 78624 77250
<< metal2 >>
rect 25536 79200 25648 80000
rect 30240 79200 30352 80000
rect 34272 79200 34384 80000
rect 34944 79200 35056 80000
rect 35616 79200 35728 80000
rect 47040 79200 47152 80000
rect 49728 79200 49840 80000
rect 50400 79200 50512 80000
rect 56448 79200 56560 80000
rect 57792 79200 57904 80000
rect 58464 79200 58576 80000
rect 59136 79200 59248 80000
rect 59808 79200 59920 80000
rect 60480 79200 60592 80000
rect 28224 0 28336 800
rect 34944 0 35056 800
rect 38304 0 38416 800
rect 48384 0 48496 800
rect 49728 0 49840 800
rect 59136 0 59248 800
rect 62496 0 62608 800
rect 63168 0 63280 800
rect 67200 0 67312 800
<< obsm2 >>
rect 4476 79140 25476 79200
rect 25708 79140 30180 79200
rect 30412 79140 34212 79200
rect 34444 79140 34884 79200
rect 35116 79140 35556 79200
rect 35788 79140 46980 79200
rect 47212 79140 49668 79200
rect 49900 79140 50340 79200
rect 50572 79140 56388 79200
rect 56620 79140 57732 79200
rect 57964 79140 58404 79200
rect 58636 79140 59076 79200
rect 59308 79140 59748 79200
rect 59980 79140 60420 79200
rect 60652 79140 78484 79200
rect 4476 860 78484 79140
rect 4476 800 28164 860
rect 28396 800 34884 860
rect 35116 800 38244 860
rect 38476 800 48324 860
rect 48556 800 49668 860
rect 49900 800 59076 860
rect 59308 800 62436 860
rect 62668 800 63108 860
rect 63340 800 67140 860
rect 67372 800 78484 860
<< metal3 >>
rect 79200 64512 80000 64624
rect 79200 60480 80000 60592
rect 79200 59808 80000 59920
rect 79200 57792 80000 57904
rect 79200 49728 80000 49840
rect 79200 47712 80000 47824
rect 79200 47040 80000 47152
rect 79200 46368 80000 46480
rect 79200 45696 80000 45808
rect 79200 45024 80000 45136
rect 79200 43008 80000 43120
rect 79200 42336 80000 42448
rect 79200 40992 80000 41104
rect 79200 40320 80000 40432
rect 79200 37632 80000 37744
rect 79200 29568 80000 29680
rect 79200 28896 80000 29008
rect 79200 28224 80000 28336
rect 79200 26880 80000 26992
rect 79200 19488 80000 19600
rect 79200 18816 80000 18928
rect 79200 16800 80000 16912
rect 79200 16128 80000 16240
rect 79200 15456 80000 15568
<< obsm3 >>
rect 4466 64684 79268 76860
rect 4466 64452 79140 64684
rect 4466 60652 79268 64452
rect 4466 60420 79140 60652
rect 4466 59980 79268 60420
rect 4466 59748 79140 59980
rect 4466 57964 79268 59748
rect 4466 57732 79140 57964
rect 4466 49900 79268 57732
rect 4466 49668 79140 49900
rect 4466 47884 79268 49668
rect 4466 47652 79140 47884
rect 4466 47212 79268 47652
rect 4466 46980 79140 47212
rect 4466 46540 79268 46980
rect 4466 46308 79140 46540
rect 4466 45868 79268 46308
rect 4466 45636 79140 45868
rect 4466 45196 79268 45636
rect 4466 44964 79140 45196
rect 4466 43180 79268 44964
rect 4466 42948 79140 43180
rect 4466 42508 79268 42948
rect 4466 42276 79140 42508
rect 4466 41164 79268 42276
rect 4466 40932 79140 41164
rect 4466 40492 79268 40932
rect 4466 40260 79140 40492
rect 4466 37804 79268 40260
rect 4466 37572 79140 37804
rect 4466 29740 79268 37572
rect 4466 29508 79140 29740
rect 4466 29068 79268 29508
rect 4466 28836 79140 29068
rect 4466 28396 79268 28836
rect 4466 28164 79140 28396
rect 4466 27052 79268 28164
rect 4466 26820 79140 27052
rect 4466 19660 79268 26820
rect 4466 19428 79140 19660
rect 4466 18988 79268 19428
rect 4466 18756 79140 18988
rect 4466 16972 79268 18756
rect 4466 16740 79140 16972
rect 4466 16300 79268 16740
rect 4466 16068 79140 16300
rect 4466 15628 79268 16068
rect 4466 15396 79140 15628
rect 4466 3108 79268 15396
<< metal4 >>
rect 4448 3076 4768 76892
rect 19808 3076 20128 76892
rect 35168 3076 35488 76892
rect 50528 3076 50848 76892
rect 65888 3076 66208 76892
<< labels >>
rlabel metal2 s 28224 0 28336 800 6 clk
port 1 nsew signal input
rlabel metal3 s 79200 40992 80000 41104 6 clk_s
port 2 nsew signal output
rlabel metal3 s 79200 47040 80000 47152 6 dir
port 3 nsew signal input
rlabel metal3 s 79200 45696 80000 45808 6 enable
port 4 nsew signal input
rlabel metal3 s 79200 26880 80000 26992 6 io_oeb[0]
port 5 nsew signal output
rlabel metal2 s 48384 0 48496 800 6 io_oeb[10]
port 6 nsew signal output
rlabel metal2 s 62496 0 62608 800 6 io_oeb[11]
port 7 nsew signal output
rlabel metal3 s 79200 49728 80000 49840 6 io_oeb[12]
port 8 nsew signal output
rlabel metal2 s 59136 79200 59248 80000 6 io_oeb[13]
port 9 nsew signal output
rlabel metal2 s 50400 79200 50512 80000 6 io_oeb[14]
port 10 nsew signal output
rlabel metal3 s 79200 28896 80000 29008 6 io_oeb[15]
port 11 nsew signal output
rlabel metal2 s 67200 0 67312 800 6 io_oeb[16]
port 12 nsew signal output
rlabel metal3 s 79200 16800 80000 16912 6 io_oeb[17]
port 13 nsew signal output
rlabel metal2 s 38304 0 38416 800 6 io_oeb[18]
port 14 nsew signal output
rlabel metal3 s 79200 43008 80000 43120 6 io_oeb[19]
port 15 nsew signal output
rlabel metal3 s 79200 29568 80000 29680 6 io_oeb[1]
port 16 nsew signal output
rlabel metal2 s 25536 79200 25648 80000 6 io_oeb[20]
port 17 nsew signal output
rlabel metal2 s 30240 79200 30352 80000 6 io_oeb[21]
port 18 nsew signal output
rlabel metal2 s 34272 79200 34384 80000 6 io_oeb[22]
port 19 nsew signal output
rlabel metal2 s 58464 79200 58576 80000 6 io_oeb[23]
port 20 nsew signal output
rlabel metal3 s 79200 57792 80000 57904 6 io_oeb[24]
port 21 nsew signal output
rlabel metal3 s 79200 16128 80000 16240 6 io_oeb[25]
port 22 nsew signal output
rlabel metal3 s 79200 19488 80000 19600 6 io_oeb[26]
port 23 nsew signal output
rlabel metal3 s 79200 64512 80000 64624 6 io_oeb[27]
port 24 nsew signal output
rlabel metal3 s 79200 28224 80000 28336 6 io_oeb[28]
port 25 nsew signal output
rlabel metal3 s 79200 46368 80000 46480 6 io_oeb[29]
port 26 nsew signal output
rlabel metal2 s 56448 79200 56560 80000 6 io_oeb[2]
port 27 nsew signal output
rlabel metal2 s 63168 0 63280 800 6 io_oeb[30]
port 28 nsew signal output
rlabel metal2 s 60480 79200 60592 80000 6 io_oeb[31]
port 29 nsew signal output
rlabel metal3 s 79200 59808 80000 59920 6 io_oeb[32]
port 30 nsew signal output
rlabel metal2 s 34944 0 35056 800 6 io_oeb[33]
port 31 nsew signal output
rlabel metal2 s 59136 0 59248 800 6 io_oeb[34]
port 32 nsew signal output
rlabel metal2 s 49728 79200 49840 80000 6 io_oeb[35]
port 33 nsew signal output
rlabel metal2 s 59808 79200 59920 80000 6 io_oeb[36]
port 34 nsew signal output
rlabel metal2 s 49728 0 49840 800 6 io_oeb[37]
port 35 nsew signal output
rlabel metal2 s 35616 79200 35728 80000 6 io_oeb[3]
port 36 nsew signal output
rlabel metal2 s 34944 79200 35056 80000 6 io_oeb[4]
port 37 nsew signal output
rlabel metal3 s 79200 60480 80000 60592 6 io_oeb[5]
port 38 nsew signal output
rlabel metal3 s 79200 18816 80000 18928 6 io_oeb[6]
port 39 nsew signal output
rlabel metal3 s 79200 15456 80000 15568 6 io_oeb[7]
port 40 nsew signal output
rlabel metal2 s 57792 79200 57904 80000 6 io_oeb[8]
port 41 nsew signal output
rlabel metal3 s 79200 37632 80000 37744 6 io_oeb[9]
port 42 nsew signal output
rlabel metal3 s 79200 40320 80000 40432 6 rst
port 43 nsew signal input
rlabel metal3 s 79200 42336 80000 42448 6 salida[0]
port 44 nsew signal output
rlabel metal3 s 79200 45024 80000 45136 6 salida[1]
port 45 nsew signal output
rlabel metal2 s 47040 79200 47152 80000 6 salida[2]
port 46 nsew signal output
rlabel metal3 s 79200 47712 80000 47824 6 salida[3]
port 47 nsew signal output
rlabel metal4 s 4448 3076 4768 76892 6 vdd
port 48 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 76892 6 vdd
port 48 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 76892 6 vdd
port 48 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 76892 6 vss
port 49 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 76892 6 vss
port 49 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 939938
string GDS_FILE /home/gf180mcu/caravel_user_project/openlane/control_system/runs/23_12_09_10_12/results/signoff/control_system.magic.gds
string GDS_START 179464
<< end >>

