VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO control_system
  CLASS BLOCK ;
  FOREIGN control_system ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END clk
  PIN clk_s
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 204.960 400.000 205.520 ;
    END
  END clk_s
  PIN dir
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 235.200 400.000 235.760 ;
    END
  END dir
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 228.480 400.000 229.040 ;
    END
  END enable
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 134.400 400.000 134.960 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 0.000 242.480 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 0.000 313.040 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 248.640 400.000 249.200 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 396.000 296.240 400.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 396.000 252.560 400.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 144.480 400.000 145.040 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 0.000 336.560 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 84.000 400.000 84.560 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 215.040 400.000 215.600 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 147.840 400.000 148.400 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 396.000 128.240 400.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 396.000 151.760 400.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 396.000 171.920 400.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 396.000 292.880 400.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 288.960 400.000 289.520 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 80.640 400.000 81.200 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 97.440 400.000 98.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 322.560 400.000 323.120 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 141.120 400.000 141.680 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 231.840 400.000 232.400 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 396.000 282.800 400.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 0.000 316.400 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 396.000 302.960 400.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 299.040 400.000 299.600 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 0.000 175.280 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 0.000 296.240 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 396.000 249.200 400.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 396.000 299.600 400.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 0.000 249.200 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 396.000 178.640 400.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 396.000 175.280 400.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 302.400 400.000 302.960 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 94.080 400.000 94.640 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 77.280 400.000 77.840 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 396.000 289.520 400.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 188.160 400.000 188.720 ;
    END
  END io_oeb[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 201.600 400.000 202.160 ;
    END
  END rst
  PIN salida[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 211.680 400.000 212.240 ;
    END
  END salida[0]
  PIN salida[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 225.120 400.000 225.680 ;
    END
  END salida[1]
  PIN salida[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 396.000 235.760 400.000 ;
    END
  END salida[2]
  PIN salida[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 396.000 238.560 400.000 239.120 ;
    END
  END salida[3]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 384.460 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 384.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 384.460 ;
    END
  END vss
  OBS
      LAYER Pwell ;
        RECT 6.290 382.400 393.550 384.590 ;
      LAYER Nwell ;
        RECT 6.290 378.080 393.550 382.400 ;
      LAYER Pwell ;
        RECT 6.290 374.560 393.550 378.080 ;
      LAYER Nwell ;
        RECT 6.290 370.240 393.550 374.560 ;
      LAYER Pwell ;
        RECT 6.290 366.720 393.550 370.240 ;
      LAYER Nwell ;
        RECT 6.290 362.400 393.550 366.720 ;
      LAYER Pwell ;
        RECT 6.290 358.880 393.550 362.400 ;
      LAYER Nwell ;
        RECT 6.290 354.560 393.550 358.880 ;
      LAYER Pwell ;
        RECT 6.290 351.040 393.550 354.560 ;
      LAYER Nwell ;
        RECT 6.290 346.720 393.550 351.040 ;
      LAYER Pwell ;
        RECT 6.290 343.200 393.550 346.720 ;
      LAYER Nwell ;
        RECT 6.290 338.880 393.550 343.200 ;
      LAYER Pwell ;
        RECT 6.290 335.360 393.550 338.880 ;
      LAYER Nwell ;
        RECT 6.290 331.040 393.550 335.360 ;
      LAYER Pwell ;
        RECT 6.290 327.520 393.550 331.040 ;
      LAYER Nwell ;
        RECT 6.290 323.200 393.550 327.520 ;
      LAYER Pwell ;
        RECT 6.290 319.680 393.550 323.200 ;
      LAYER Nwell ;
        RECT 6.290 315.360 393.550 319.680 ;
      LAYER Pwell ;
        RECT 6.290 311.840 393.550 315.360 ;
      LAYER Nwell ;
        RECT 6.290 307.520 393.550 311.840 ;
      LAYER Pwell ;
        RECT 6.290 304.000 393.550 307.520 ;
      LAYER Nwell ;
        RECT 6.290 299.680 393.550 304.000 ;
      LAYER Pwell ;
        RECT 6.290 296.160 393.550 299.680 ;
      LAYER Nwell ;
        RECT 6.290 291.840 393.550 296.160 ;
      LAYER Pwell ;
        RECT 6.290 288.320 393.550 291.840 ;
      LAYER Nwell ;
        RECT 6.290 284.000 393.550 288.320 ;
      LAYER Pwell ;
        RECT 6.290 280.480 393.550 284.000 ;
      LAYER Nwell ;
        RECT 6.290 276.160 393.550 280.480 ;
      LAYER Pwell ;
        RECT 6.290 272.640 393.550 276.160 ;
      LAYER Nwell ;
        RECT 6.290 268.320 393.550 272.640 ;
      LAYER Pwell ;
        RECT 6.290 264.800 393.550 268.320 ;
      LAYER Nwell ;
        RECT 6.290 260.480 393.550 264.800 ;
      LAYER Pwell ;
        RECT 6.290 256.960 393.550 260.480 ;
      LAYER Nwell ;
        RECT 6.290 252.640 393.550 256.960 ;
      LAYER Pwell ;
        RECT 6.290 249.120 393.550 252.640 ;
      LAYER Nwell ;
        RECT 6.290 244.925 393.550 249.120 ;
        RECT 6.290 244.800 228.305 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 393.550 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 257.985 241.280 ;
        RECT 6.290 237.085 393.550 241.155 ;
        RECT 6.290 236.960 168.945 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 393.550 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 145.985 233.440 ;
        RECT 6.290 229.245 393.550 233.315 ;
        RECT 6.290 229.120 149.905 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 393.550 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 151.630 225.600 ;
        RECT 6.290 221.405 393.550 225.475 ;
        RECT 6.290 221.280 210.945 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 393.550 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 190.880 217.760 ;
        RECT 6.290 213.565 393.550 217.635 ;
        RECT 6.290 213.440 149.905 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 393.550 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 143.745 209.920 ;
        RECT 6.290 205.725 393.550 209.795 ;
        RECT 6.290 205.600 205.000 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 393.550 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 184.280 202.080 ;
        RECT 6.290 197.885 393.550 201.955 ;
        RECT 6.290 197.760 206.120 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 393.550 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 152.145 194.240 ;
        RECT 6.290 190.045 393.550 194.115 ;
        RECT 6.290 189.920 154.430 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 393.550 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 148.785 186.400 ;
        RECT 6.290 182.205 393.550 186.275 ;
        RECT 6.290 182.080 171.745 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 393.550 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 216.545 178.560 ;
        RECT 6.290 174.365 393.550 178.435 ;
        RECT 6.290 174.240 149.905 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 393.550 174.240 ;
      LAYER Nwell ;
        RECT 6.290 166.400 393.550 170.720 ;
      LAYER Pwell ;
        RECT 6.290 162.880 393.550 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 151.630 162.880 ;
        RECT 6.290 158.685 393.550 162.755 ;
        RECT 6.290 158.560 166.920 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 393.550 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 144.305 155.040 ;
        RECT 6.290 150.720 393.550 154.915 ;
      LAYER Pwell ;
        RECT 6.290 147.200 393.550 150.720 ;
      LAYER Nwell ;
        RECT 6.290 143.005 393.550 147.200 ;
        RECT 6.290 142.880 151.025 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 393.550 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 157.790 139.360 ;
        RECT 6.290 135.040 393.550 139.235 ;
      LAYER Pwell ;
        RECT 6.290 131.520 393.550 135.040 ;
      LAYER Nwell ;
        RECT 6.290 127.200 393.550 131.520 ;
      LAYER Pwell ;
        RECT 6.290 123.680 393.550 127.200 ;
      LAYER Nwell ;
        RECT 6.290 119.360 393.550 123.680 ;
      LAYER Pwell ;
        RECT 6.290 115.840 393.550 119.360 ;
      LAYER Nwell ;
        RECT 6.290 111.520 393.550 115.840 ;
      LAYER Pwell ;
        RECT 6.290 108.000 393.550 111.520 ;
      LAYER Nwell ;
        RECT 6.290 103.680 393.550 108.000 ;
      LAYER Pwell ;
        RECT 6.290 100.160 393.550 103.680 ;
      LAYER Nwell ;
        RECT 6.290 95.840 393.550 100.160 ;
      LAYER Pwell ;
        RECT 6.290 92.320 393.550 95.840 ;
      LAYER Nwell ;
        RECT 6.290 88.000 393.550 92.320 ;
      LAYER Pwell ;
        RECT 6.290 84.480 393.550 88.000 ;
      LAYER Nwell ;
        RECT 6.290 80.160 393.550 84.480 ;
      LAYER Pwell ;
        RECT 6.290 76.640 393.550 80.160 ;
      LAYER Nwell ;
        RECT 6.290 72.320 393.550 76.640 ;
      LAYER Pwell ;
        RECT 6.290 68.800 393.550 72.320 ;
      LAYER Nwell ;
        RECT 6.290 64.480 393.550 68.800 ;
      LAYER Pwell ;
        RECT 6.290 60.960 393.550 64.480 ;
      LAYER Nwell ;
        RECT 6.290 56.640 393.550 60.960 ;
      LAYER Pwell ;
        RECT 6.290 53.120 393.550 56.640 ;
      LAYER Nwell ;
        RECT 6.290 48.800 393.550 53.120 ;
      LAYER Pwell ;
        RECT 6.290 45.280 393.550 48.800 ;
      LAYER Nwell ;
        RECT 6.290 40.960 393.550 45.280 ;
      LAYER Pwell ;
        RECT 6.290 37.440 393.550 40.960 ;
      LAYER Nwell ;
        RECT 6.290 33.120 393.550 37.440 ;
      LAYER Pwell ;
        RECT 6.290 29.600 393.550 33.120 ;
      LAYER Nwell ;
        RECT 6.290 25.280 393.550 29.600 ;
      LAYER Pwell ;
        RECT 6.290 21.760 393.550 25.280 ;
      LAYER Nwell ;
        RECT 6.290 17.440 393.550 21.760 ;
      LAYER Pwell ;
        RECT 6.290 15.250 393.550 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 393.120 386.250 ;
      LAYER Metal2 ;
        RECT 22.380 395.700 127.380 396.000 ;
        RECT 128.540 395.700 150.900 396.000 ;
        RECT 152.060 395.700 171.060 396.000 ;
        RECT 172.220 395.700 174.420 396.000 ;
        RECT 175.580 395.700 177.780 396.000 ;
        RECT 178.940 395.700 234.900 396.000 ;
        RECT 236.060 395.700 248.340 396.000 ;
        RECT 249.500 395.700 251.700 396.000 ;
        RECT 252.860 395.700 281.940 396.000 ;
        RECT 283.100 395.700 288.660 396.000 ;
        RECT 289.820 395.700 292.020 396.000 ;
        RECT 293.180 395.700 295.380 396.000 ;
        RECT 296.540 395.700 298.740 396.000 ;
        RECT 299.900 395.700 302.100 396.000 ;
        RECT 303.260 395.700 392.420 396.000 ;
        RECT 22.380 4.300 392.420 395.700 ;
        RECT 22.380 4.000 140.820 4.300 ;
        RECT 141.980 4.000 174.420 4.300 ;
        RECT 175.580 4.000 191.220 4.300 ;
        RECT 192.380 4.000 241.620 4.300 ;
        RECT 242.780 4.000 248.340 4.300 ;
        RECT 249.500 4.000 295.380 4.300 ;
        RECT 296.540 4.000 312.180 4.300 ;
        RECT 313.340 4.000 315.540 4.300 ;
        RECT 316.700 4.000 335.700 4.300 ;
        RECT 336.860 4.000 392.420 4.300 ;
      LAYER Metal3 ;
        RECT 22.330 323.420 396.340 384.300 ;
        RECT 22.330 322.260 395.700 323.420 ;
        RECT 22.330 303.260 396.340 322.260 ;
        RECT 22.330 302.100 395.700 303.260 ;
        RECT 22.330 299.900 396.340 302.100 ;
        RECT 22.330 298.740 395.700 299.900 ;
        RECT 22.330 289.820 396.340 298.740 ;
        RECT 22.330 288.660 395.700 289.820 ;
        RECT 22.330 249.500 396.340 288.660 ;
        RECT 22.330 248.340 395.700 249.500 ;
        RECT 22.330 239.420 396.340 248.340 ;
        RECT 22.330 238.260 395.700 239.420 ;
        RECT 22.330 236.060 396.340 238.260 ;
        RECT 22.330 234.900 395.700 236.060 ;
        RECT 22.330 232.700 396.340 234.900 ;
        RECT 22.330 231.540 395.700 232.700 ;
        RECT 22.330 229.340 396.340 231.540 ;
        RECT 22.330 228.180 395.700 229.340 ;
        RECT 22.330 225.980 396.340 228.180 ;
        RECT 22.330 224.820 395.700 225.980 ;
        RECT 22.330 215.900 396.340 224.820 ;
        RECT 22.330 214.740 395.700 215.900 ;
        RECT 22.330 212.540 396.340 214.740 ;
        RECT 22.330 211.380 395.700 212.540 ;
        RECT 22.330 205.820 396.340 211.380 ;
        RECT 22.330 204.660 395.700 205.820 ;
        RECT 22.330 202.460 396.340 204.660 ;
        RECT 22.330 201.300 395.700 202.460 ;
        RECT 22.330 189.020 396.340 201.300 ;
        RECT 22.330 187.860 395.700 189.020 ;
        RECT 22.330 148.700 396.340 187.860 ;
        RECT 22.330 147.540 395.700 148.700 ;
        RECT 22.330 145.340 396.340 147.540 ;
        RECT 22.330 144.180 395.700 145.340 ;
        RECT 22.330 141.980 396.340 144.180 ;
        RECT 22.330 140.820 395.700 141.980 ;
        RECT 22.330 135.260 396.340 140.820 ;
        RECT 22.330 134.100 395.700 135.260 ;
        RECT 22.330 98.300 396.340 134.100 ;
        RECT 22.330 97.140 395.700 98.300 ;
        RECT 22.330 94.940 396.340 97.140 ;
        RECT 22.330 93.780 395.700 94.940 ;
        RECT 22.330 84.860 396.340 93.780 ;
        RECT 22.330 83.700 395.700 84.860 ;
        RECT 22.330 81.500 396.340 83.700 ;
        RECT 22.330 80.340 395.700 81.500 ;
        RECT 22.330 78.140 396.340 80.340 ;
        RECT 22.330 76.980 395.700 78.140 ;
        RECT 22.330 15.540 396.340 76.980 ;
  END
END control_system
END LIBRARY

