// This is the unpowered netlist.
module control_system (clk,
    clk_s,
    dir,
    enable,
    rst,
    io_oeb,
    salida);
 input clk;
 output clk_s;
 input dir;
 input enable;
 input rst;
 output [37:0] io_oeb;
 output [3:0] salida;

 wire net44;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net45;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net46;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net13;
 wire net14;
 wire net15;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire \count[0] ;
 wire \count[10] ;
 wire \count[11] ;
 wire \count[12] ;
 wire \count[13] ;
 wire \count[14] ;
 wire \count[15] ;
 wire \count[16] ;
 wire \count[17] ;
 wire \count[18] ;
 wire \count[19] ;
 wire \count[1] ;
 wire \count[20] ;
 wire \count[21] ;
 wire \count[22] ;
 wire \count[23] ;
 wire \count[24] ;
 wire \count[25] ;
 wire \count[26] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \count[5] ;
 wire \count[6] ;
 wire \count[7] ;
 wire \count[8] ;
 wire \count[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state_next[0] ;
 wire \state_next[1] ;
 wire \state_next[2] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout11_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(dir));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(enable));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output4_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output5_I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_292 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _154_ (.I(\count[0] ),
    .Z(_135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _155_ (.I(\count[22] ),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _156_ (.A1(\count[20] ),
    .A2(\count[21] ),
    .A3(_136_),
    .A4(\count[23] ),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _157_ (.A1(\count[16] ),
    .A2(\count[17] ),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _158_ (.A1(\count[18] ),
    .A2(\count[19] ),
    .A3(_137_),
    .A4(_138_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _159_ (.A1(\count[24] ),
    .A2(\count[25] ),
    .A3(\count[26] ),
    .A4(_139_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _160_ (.A1(\count[2] ),
    .A2(\count[3] ),
    .A3(\count[4] ),
    .A4(\count[5] ),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _161_ (.A1(\count[8] ),
    .A2(\count[9] ),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _162_ (.A1(_135_),
    .A2(\count[1] ),
    .A3(_142_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _163_ (.I(\count[15] ),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _164_ (.A1(\count[14] ),
    .A2(_144_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _165_ (.I(\count[7] ),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _166_ (.I(\count[10] ),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _167_ (.A1(\count[6] ),
    .A2(_146_),
    .A3(_147_),
    .A4(\count[11] ),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _168_ (.A1(\count[12] ),
    .A2(\count[13] ),
    .A3(_145_),
    .A4(_148_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _169_ (.A1(_140_),
    .A2(_141_),
    .A3(_143_),
    .A4(_149_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _170_ (.A1(net3),
    .A2(_150_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _171_ (.I(_151_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _172_ (.I(_152_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _173_ (.A1(_135_),
    .A2(_153_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _174_ (.A1(_135_),
    .A2(\count[1] ),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _175_ (.I(_151_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _176_ (.I(_039_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _177_ (.A1(_135_),
    .A2(\count[1] ),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _178_ (.A1(_038_),
    .A2(_040_),
    .A3(_041_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _179_ (.A1(\count[2] ),
    .A2(_041_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _180_ (.A1(_153_),
    .A2(_042_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _181_ (.I(_039_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _182_ (.A1(\count[0] ),
    .A2(\count[1] ),
    .A3(\count[2] ),
    .A4(\count[3] ),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _183_ (.I(_044_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _184_ (.A1(\count[2] ),
    .A2(_041_),
    .B(\count[3] ),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _185_ (.A1(_043_),
    .A2(_045_),
    .A3(_046_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _186_ (.A1(\count[4] ),
    .A2(_045_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _187_ (.A1(_153_),
    .A2(_047_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _188_ (.A1(\count[4] ),
    .A2(\count[5] ),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _189_ (.A1(_045_),
    .A2(_048_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _190_ (.A1(\count[4] ),
    .A2(_045_),
    .B(\count[5] ),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _191_ (.A1(_043_),
    .A2(_049_),
    .A3(_050_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _192_ (.A1(\count[6] ),
    .A2(_049_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _193_ (.A1(\count[6] ),
    .A2(_049_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _194_ (.A1(_043_),
    .A2(_051_),
    .A3(_052_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _195_ (.I(_039_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _196_ (.A1(_146_),
    .A2(_051_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _197_ (.A1(_053_),
    .A2(_054_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _198_ (.A1(\count[6] ),
    .A2(\count[7] ),
    .A3(_044_),
    .A4(_048_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _199_ (.A1(\count[8] ),
    .A2(_055_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _200_ (.A1(_053_),
    .A2(_056_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _201_ (.I(\count[9] ),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _202_ (.A1(\count[7] ),
    .A2(\count[8] ),
    .A3(_051_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _203_ (.A1(_142_),
    .A2(_055_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _204_ (.A1(_057_),
    .A2(_058_),
    .B(_059_),
    .C(_043_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _205_ (.I(_039_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _206_ (.A1(\count[10] ),
    .A2(_059_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _207_ (.A1(_147_),
    .A2(_142_),
    .A3(_055_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _208_ (.A1(_060_),
    .A2(_061_),
    .A3(_062_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _209_ (.I(\count[11] ),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _210_ (.A1(_147_),
    .A2(_063_),
    .A3(_142_),
    .A4(_055_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _211_ (.I(_064_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _212_ (.A1(\count[11] ),
    .A2(_062_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _213_ (.A1(_060_),
    .A2(_065_),
    .A3(_066_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _214_ (.A1(\count[12] ),
    .A2(_065_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _215_ (.A1(_053_),
    .A2(_067_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _216_ (.A1(\count[12] ),
    .A2(_065_),
    .B(\count[13] ),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _217_ (.A1(\count[12] ),
    .A2(\count[13] ),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _218_ (.A1(_065_),
    .A2(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _219_ (.A1(_060_),
    .A2(_068_),
    .A3(_070_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _220_ (.A1(\count[14] ),
    .A2(_070_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _221_ (.A1(_053_),
    .A2(_071_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _222_ (.A1(\count[14] ),
    .A2(\count[15] ),
    .A3(_064_),
    .A4(_069_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _223_ (.I(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _224_ (.A1(\count[14] ),
    .A2(_070_),
    .B(\count[15] ),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _225_ (.A1(_060_),
    .A2(_073_),
    .A3(_074_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _226_ (.A1(\count[16] ),
    .A2(_073_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _227_ (.A1(_040_),
    .A2(_075_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _228_ (.I(_151_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _229_ (.A1(\count[16] ),
    .A2(_073_),
    .B(\count[17] ),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _230_ (.A1(\count[16] ),
    .A2(\count[17] ),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _231_ (.A1(_073_),
    .A2(_078_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _232_ (.A1(_076_),
    .A2(_077_),
    .A3(_079_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _233_ (.A1(\count[18] ),
    .A2(_079_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _234_ (.A1(\count[18] ),
    .A2(_079_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _235_ (.A1(_076_),
    .A2(_080_),
    .A3(_081_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _236_ (.A1(\count[18] ),
    .A2(\count[19] ),
    .A3(_072_),
    .A4(_078_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _237_ (.I(_082_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _238_ (.A1(\count[19] ),
    .A2(_080_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _239_ (.A1(_076_),
    .A2(_083_),
    .A3(_084_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _240_ (.A1(\count[20] ),
    .A2(_083_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _241_ (.A1(_040_),
    .A2(_085_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _242_ (.A1(\count[20] ),
    .A2(_083_),
    .B(\count[21] ),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _243_ (.A1(\count[20] ),
    .A2(\count[21] ),
    .Z(_087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _244_ (.A1(_082_),
    .A2(_087_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _245_ (.A1(_076_),
    .A2(_086_),
    .A3(_088_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _246_ (.A1(_136_),
    .A2(_088_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _247_ (.A1(_040_),
    .A2(_089_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _248_ (.A1(\count[22] ),
    .A2(\count[23] ),
    .A3(_083_),
    .A4(_087_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _249_ (.A1(\count[22] ),
    .A2(_088_),
    .B(\count[23] ),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _250_ (.A1(_152_),
    .A2(_090_),
    .A3(_091_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _251_ (.I(\count[24] ),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _252_ (.A1(\count[22] ),
    .A2(\count[23] ),
    .A3(_082_),
    .A4(_087_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _253_ (.A1(_092_),
    .A2(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _254_ (.A1(\count[24] ),
    .A2(_090_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _255_ (.A1(_152_),
    .A2(_094_),
    .A3(_095_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _256_ (.I(\count[25] ),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _257_ (.A1(_092_),
    .A2(_096_),
    .A3(_093_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _258_ (.A1(\count[24] ),
    .A2(_090_),
    .B(\count[25] ),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _259_ (.A1(_152_),
    .A2(_097_),
    .A3(_098_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _260_ (.A1(_092_),
    .A2(_096_),
    .A3(_093_),
    .B(\count[26] ),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _261_ (.A1(_092_),
    .A2(_096_),
    .A3(\count[26] ),
    .A4(_093_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _262_ (.A1(_099_),
    .A2(_100_),
    .B(_153_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _263_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _264_ (.A1(\state[2] ),
    .A2(_101_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _265_ (.A1(\state[2] ),
    .A2(_101_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _266_ (.I(\state[0] ),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _267_ (.I(\state[2] ),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _268_ (.A1(\state[1] ),
    .A2(_104_),
    .A3(_105_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _269_ (.A1(_103_),
    .A2(_106_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _270_ (.A1(_102_),
    .A2(_107_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _271_ (.I(_108_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _272_ (.A1(net5),
    .A2(_109_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _273_ (.A1(\state[1] ),
    .A2(\state[2] ),
    .A3(_101_),
    .B(_110_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _274_ (.A1(\state[1] ),
    .A2(_105_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _275_ (.A1(net6),
    .A2(_109_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _276_ (.A1(_104_),
    .A2(_111_),
    .B(_112_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _277_ (.I(_108_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _278_ (.A1(net7),
    .A2(_113_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _279_ (.A1(_106_),
    .A2(_114_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _280_ (.I(net8),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _281_ (.I(_103_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _282_ (.A1(_115_),
    .A2(_116_),
    .B(_102_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _283_ (.A1(net2),
    .A2(_104_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _284_ (.A1(\state_next[0] ),
    .A2(_109_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _285_ (.A1(_113_),
    .A2(_117_),
    .B(_118_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _286_ (.I(\state_next[1] ),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _287_ (.I(net2),
    .Z(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _288_ (.I(_106_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _289_ (.A1(net1),
    .A2(net2),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _290_ (.A1(_120_),
    .A2(_121_),
    .B(_107_),
    .C(_122_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _291_ (.A1(net1),
    .A2(_120_),
    .A3(_116_),
    .A4(_111_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _292_ (.I(net1),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _293_ (.A1(_125_),
    .A2(_120_),
    .B(_104_),
    .C(_111_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _294_ (.A1(_108_),
    .A2(_124_),
    .A3(_126_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _295_ (.A1(_119_),
    .A2(_113_),
    .B1(_123_),
    .B2(_127_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _296_ (.I(\state_next[2] ),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _297_ (.A1(_125_),
    .A2(net2),
    .A3(_116_),
    .A4(_111_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _298_ (.A1(_120_),
    .A2(_116_),
    .B1(_106_),
    .B2(_122_),
    .C(_129_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _299_ (.A1(_109_),
    .A2(_130_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _300_ (.A1(_128_),
    .A2(_113_),
    .B(_131_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _301_ (.I(net3),
    .Z(_132_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _302_ (.A1(_132_),
    .A2(\state_next[0] ),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _303_ (.I(_133_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _304_ (.A1(_132_),
    .A2(_119_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _305_ (.A1(_132_),
    .A2(_128_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _306_ (.A1(net9),
    .A2(_150_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _307_ (.A1(_132_),
    .A2(_134_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _308_ (.D(_000_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _309_ (.D(_001_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _310_ (.D(_002_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _311_ (.D(_003_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _312_ (.D(_004_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _313_ (.D(_005_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _314_ (.D(_006_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _315_ (.D(_007_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _316_ (.D(_008_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _317_ (.D(_009_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\count[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _318_ (.D(_010_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _319_ (.D(_011_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _320_ (.D(_012_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _321_ (.D(_013_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _322_ (.D(_014_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _323_ (.D(_015_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _324_ (.D(_016_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\count[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _325_ (.D(_017_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _326_ (.D(_018_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _327_ (.D(_019_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _328_ (.D(_020_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _329_ (.D(_021_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _330_ (.D(_022_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\count[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _331_ (.D(_023_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _332_ (.D(_024_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _333_ (.D(_025_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _334_ (.D(_026_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\count[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _335_ (.D(_027_),
    .CLK(net10),
    .Q(net5));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _336_ (.D(_028_),
    .CLK(net10),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _337_ (.D(_029_),
    .CLK(net9),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _338_ (.D(_030_),
    .CLK(net10),
    .Q(net8));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _339_ (.D(_031_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state_next[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _340_ (.D(_032_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state_next[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _341_ (.D(_033_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state_next[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _342_ (.D(_034_),
    .CLK(net10),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _343_ (.D(_035_),
    .CLK(net9),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _344_ (.D(_036_),
    .CLK(net9),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _345_ (.D(_037_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_13 (.ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_14 (.ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_15 (.ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_16 (.ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_17 (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_18 (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_19 (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_20 (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_21 (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel control_system_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_44 (.Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_45 (.Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_46 (.Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_47 (.Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_48 (.Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_49 (.Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__tieh control_system_50 (.Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout10 (.I(net11),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout11 (.I(net12),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout12 (.I(net4),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout9 (.I(net11),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(dir),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(rst),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output4 (.I(net12),
    .Z(clk_s));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output5 (.I(net5),
    .Z(salida[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output6 (.I(net6),
    .Z(salida[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output7 (.I(net7),
    .Z(salida[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output8 (.I(net8),
    .Z(salida[3]));
 assign io_oeb[0] = net44;
 assign io_oeb[10] = net16;
 assign io_oeb[11] = net17;
 assign io_oeb[12] = net18;
 assign io_oeb[13] = net19;
 assign io_oeb[14] = net20;
 assign io_oeb[15] = net21;
 assign io_oeb[16] = net22;
 assign io_oeb[17] = net23;
 assign io_oeb[18] = net24;
 assign io_oeb[19] = net25;
 assign io_oeb[1] = net45;
 assign io_oeb[20] = net26;
 assign io_oeb[21] = net27;
 assign io_oeb[22] = net28;
 assign io_oeb[23] = net29;
 assign io_oeb[24] = net30;
 assign io_oeb[25] = net31;
 assign io_oeb[26] = net32;
 assign io_oeb[27] = net33;
 assign io_oeb[28] = net34;
 assign io_oeb[29] = net35;
 assign io_oeb[2] = net46;
 assign io_oeb[30] = net36;
 assign io_oeb[31] = net37;
 assign io_oeb[32] = net38;
 assign io_oeb[33] = net39;
 assign io_oeb[34] = net40;
 assign io_oeb[35] = net41;
 assign io_oeb[36] = net42;
 assign io_oeb[37] = net43;
 assign io_oeb[3] = net47;
 assign io_oeb[4] = net48;
 assign io_oeb[5] = net49;
 assign io_oeb[6] = net50;
 assign io_oeb[7] = net13;
 assign io_oeb[8] = net14;
 assign io_oeb[9] = net15;
endmodule

